{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(to bottom, #fff394 0%, rgb(252,228,172) 100%)", "background-pattern":"" , "items": [ {"x": -376,"y": -2,"w": 2313,"h": 472,"type":"text","text": "","text-data": "{title}","font": "roboto condensed","color": "rgb(232,158,33)","font-size": 37, "font-style":"bold", "justification": 0 }, {"x": -368,"y": 296,"w": 2130,"h": 243,"type":"text","text": "","text-data": "{subtitle}","font": "raleway","color": "rgba(0,0,0,0.40493)","font-size": 21, "font-style":"medium", "justification": 0 }, {"x": -373,"y": 511,"w": 2239,"h": 860,"type":"image", "image":"jpg", "image-data":"/9j/4AAQSkZJRgABAQEASABIAAD/4gxYSUNDX1BST0ZJTEUAAQEAAAxITGlubwIQAABtbnRyUkdCIFhZWiAHzgACAAkABgAxAABhY3NwTVNGVAAAAABJRUMgc1JHQgAAAAAAAAAAAAAAAAAA9tYAAQAAAADTLUhQICAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABFjcHJ0AAABUAAAADNkZXNjAAABhAAAAGx3dHB0AAAB8AAAABRia3B0AAACBAAAABRyWFlaAAACGAAAABRnWFlaAAACLAAAABRiWFlaAAACQAAAABRkbW5kAAACVAAAAHBkbWRkAAACxAAAAIh2dWVkAAADTAAAAIZ2aWV3AAAD1AAAACRsdW1pAAAD+AAAABRtZWFzAAAEDAAAACR0ZWNoAAAEMAAAAAxyVFJDAAAEPAAACAxnVFJDAAAEPAAACAxiVFJDAAAEPAAACAx0ZXh0AAAAAENvcHlyaWdodCAoYykgMTk5OCBIZXdsZXR0LVBhY2thcmQgQ29tcGFueQAAZGVzYwAAAAAAAAASc1JHQiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAABJzUkdCIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAWFlaIAAAAAAAAPNRAAEAAAABFsxYWVogAAAAAAAAAAAAAAAAAAAAAFhZWiAAAAAAAABvogAAOPUAAAOQWFlaIAAAAAAAAGKZAAC3hQAAGNpYWVogAAAAAAAAJKAAAA+EAAC2z2Rlc2MAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABkZXNjAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAAAAAAAAAAAAAAAAZGVzYwAAAAAAAAAsUmVmZXJlbmNlIFZpZXdpbmcgQ29uZGl0aW9uIGluIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAALFJlZmVyZW5jZSBWaWV3aW5nIENvbmRpdGlvbiBpbiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAHZpZXcAAAAAABOk/gAUXy4AEM8UAAPtzAAEEwsAA1yeAAAAAVhZWiAAAAAAAEwJVgBQAAAAVx/nbWVhcwAAAAAAAAABAAAAAAAAAAAAAAAAAAAAAAAAAo8AAAACc2lnIAAAAABDUlQgY3VydgAAAAAAAAQAAAAABQAKAA8AFAAZAB4AIwAoAC0AMgA3ADsAQABFAEoATwBUAFkAXgBjAGgAbQByAHcAfACBAIYAiwCQAJUAmgCfAKQAqQCuALIAtwC8AMEAxgDLANAA1QDbAOAA5QDrAPAA9gD7AQEBBwENARMBGQEfASUBKwEyATgBPgFFAUwBUgFZAWABZwFuAXUBfAGDAYsBkgGaAaEBqQGxAbkBwQHJAdEB2QHhAekB8gH6AgMCDAIUAh0CJgIvAjgCQQJLAlQCXQJnAnECegKEAo4CmAKiAqwCtgLBAssC1QLgAusC9QMAAwsDFgMhAy0DOANDA08DWgNmA3IDfgOKA5YDogOuA7oDxwPTA+AD7AP5BAYEEwQgBC0EOwRIBFUEYwRxBH4EjASaBKgEtgTEBNME4QTwBP4FDQUcBSsFOgVJBVgFZwV3BYYFlgWmBbUFxQXVBeUF9gYGBhYGJwY3BkgGWQZqBnsGjAadBq8GwAbRBuMG9QcHBxkHKwc9B08HYQd0B4YHmQesB78H0gflB/gICwgfCDIIRghaCG4IggiWCKoIvgjSCOcI+wkQCSUJOglPCWQJeQmPCaQJugnPCeUJ+woRCicKPQpUCmoKgQqYCq4KxQrcCvMLCwsiCzkLUQtpC4ALmAuwC8gL4Qv5DBIMKgxDDFwMdQyODKcMwAzZDPMNDQ0mDUANWg10DY4NqQ3DDd4N+A4TDi4OSQ5kDn8Omw62DtIO7g8JDyUPQQ9eD3oPlg+zD88P7BAJECYQQxBhEH4QmxC5ENcQ9RETETERTxFtEYwRqhHJEegSBxImEkUSZBKEEqMSwxLjEwMTIxNDE2MTgxOkE8UT5RQGFCcUSRRqFIsUrRTOFPAVEhU0FVYVeBWbFb0V4BYDFiYWSRZsFo8WshbWFvoXHRdBF2UXiReuF9IX9xgbGEAYZRiKGK8Y1Rj6GSAZRRlrGZEZtxndGgQaKhpRGncanhrFGuwbFBs7G2MbihuyG9ocAhwqHFIcexyjHMwc9R0eHUcdcB2ZHcMd7B4WHkAeah6UHr4e6R8THz4faR+UH78f6iAVIEEgbCCYIMQg8CEcIUghdSGhIc4h+yInIlUigiKvIt0jCiM4I2YjlCPCI/AkHyRNJHwkqyTaJQklOCVoJZclxyX3JicmVyaHJrcm6CcYJ0kneierJ9woDSg/KHEooijUKQYpOClrKZ0p0CoCKjUqaCqbKs8rAis2K2krnSvRLAUsOSxuLKIs1y0MLUEtdi2rLeEuFi5MLoIuty7uLyQvWi+RL8cv/jA1MGwwpDDbMRIxSjGCMbox8jIqMmMymzLUMw0zRjN/M7gz8TQrNGU0njTYNRM1TTWHNcI1/TY3NnI2rjbpNyQ3YDecN9c4FDhQOIw4yDkFOUI5fzm8Ofk6Njp0OrI67zstO2s7qjvoPCc8ZTykPOM9Ij1hPaE94D4gPmA+oD7gPyE/YT+iP+JAI0BkQKZA50EpQWpBrEHuQjBCckK1QvdDOkN9Q8BEA0RHRIpEzkUSRVVFmkXeRiJGZ0arRvBHNUd7R8BIBUhLSJFI10kdSWNJqUnwSjdKfUrESwxLU0uaS+JMKkxyTLpNAk1KTZNN3E4lTm5Ot08AT0lPk0/dUCdQcVC7UQZRUFGbUeZSMVJ8UsdTE1NfU6pT9lRCVI9U21UoVXVVwlYPVlxWqVb3V0RXklfgWC9YfVjLWRpZaVm4WgdaVlqmWvVbRVuVW+VcNVyGXNZdJ114XcleGl5sXr1fD19hX7NgBWBXYKpg/GFPYaJh9WJJYpxi8GNDY5dj62RAZJRk6WU9ZZJl52Y9ZpJm6Gc9Z5Nn6Wg/aJZo7GlDaZpp8WpIap9q92tPa6dr/2xXbK9tCG1gbbluEm5rbsRvHm94b9FwK3CGcOBxOnGVcfByS3KmcwFzXXO4dBR0cHTMdSh1hXXhdj52m3b4d1Z3s3gReG54zHkqeYl553pGeqV7BHtje8J8IXyBfOF9QX2hfgF+Yn7CfyN/hH/lgEeAqIEKgWuBzYIwgpKC9INXg7qEHYSAhOOFR4Wrhg6GcobXhzuHn4gEiGmIzokziZmJ/opkisqLMIuWi/yMY4zKjTGNmI3/jmaOzo82j56QBpBukNaRP5GokhGSepLjk02TtpQglIqU9JVflcmWNJaflwqXdZfgmEyYuJkkmZCZ/JpomtWbQpuvnByciZz3nWSd0p5Anq6fHZ+Ln/qgaaDYoUehtqImopajBqN2o+akVqTHpTilqaYapoum/adup+CoUqjEqTepqaocqo+rAqt1q+msXKzQrUStuK4trqGvFq+LsACwdbDqsWCx1rJLssKzOLOutCW0nLUTtYq2AbZ5tvC3aLfguFm40blKucK6O7q1uy67p7whvJu9Fb2Pvgq+hL7/v3q/9cBwwOzBZ8Hjwl/C28NYw9TEUcTOxUvFyMZGxsPHQce/yD3IvMk6ybnKOMq3yzbLtsw1zLXNNc21zjbOts83z7jQOdC60TzRvtI/0sHTRNPG1EnUy9VO1dHWVdbY11zX4Nhk2OjZbNnx2nba+9uA3AXcit0Q3ZbeHN6i3ynfr+A24L3hROHM4lPi2+Nj4+vkc+T85YTmDeaW5x/nqegy6LzpRunQ6lvq5etw6/vshu0R7ZzuKO6070DvzPBY8OXxcvH/8ozzGfOn9DT0wvVQ9d72bfb794r4Gfio+Tj5x/pX+uf7d/wH/Jj9Kf26/kv+3P9t////2wBDAAMCAgMCAgMDAwMEAwMEBQgFBQQEBQoHBwYIDAoMDAsKCwsNDhIQDQ4RDgsLEBYQERMUFRUVDA8XGBYUGBIUFRT/2wBDAQMEBAUEBQkFBQkUDQsNFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBT/wgARCAH2BZIDAREAAhEBAxEB/8QAHAAAAwEBAQEBAQAAAAAAAAAAAAECAwQFBgcI/8QAGgEBAQEBAQEBAAAAAAAAAAAAAAECAwQFBv/aAAwDAQACEAMQAAAB/dfzf04xqyrKLLR21V2UlF07LsqnZdy9R6lWVZVhZVlXNUajsKdhoD0YUAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAATkQQZqhSkqylVmyqlUsyqVSqJlUqlUskqoRJIhCEICQAVAoQkQCFaoKUFJABAIQCAViQEAAKikJQQgRCCEAggEKgRIqUu/XPoePtGNUWlVZRWlo6tKK1LppWpVlWPWXZVlWOyrHqVY6LHY6NQp06KAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAhCggyUpCzoiYmaUqlRMsyk1MLNlVmizESoRIlmBESqsQgEAoKlBVCpAIQAJClBQAhAIBWIAEgAgoEqRWkKkgEIQCgEFKEqsRJv0noeXtPPVFJZdOrqkqrkrSrKsoepVlay7KsqyrCytR2VY6LHY6NQoK0AoAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAFkoIJVkpSVZSs5qlUsyzKlJZlnNUqlUSqJFCJpSqBJpUhAIBQUpEpYhQWoQCASAgohUCAQCsBCAEBCChUIVAkJUiCBUiBUiFahRtvHoebvPPVVSWtjqrKspbS7HVWXY9SkrUdj1mrKsdlWPUpHoWNDR6hQPRhQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAATkQQZqhSks5TKpVKpZlmaBSzKpZlJVEwlkQlUk0pQQkQhUgEACFCokSoVIBAIEQgoEoiACbAQCABBQIQhAIQSAlSCoQhCVJt0noeXrHPV1RZZVlW1ZRSUlaVZdlU7mrHqOyrKsdjsdlWOytCxoaOw0B06KAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACFCgglWaoJVE5qWZVmoUszShSqWVWapUTKhCVSSJUIIVkipCABCgESIBUQUhCQURColVCCgkVgKASCoKSghUQgEiBEoAhQE2oQjbee7zdZ56qrKKS1unZVUUlJWlWXYx6lXNajsdl2Ox2VY9SrHYWOnqGgOnRQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAQoUEGaskpLOSlmVSqVLOalUqic6lSFmysihCJWQhCETSQFQAoQCEIQgVICAVIEQKgoEAIAISAhAFqkVoIBQrAQAIBQhKhUo26zt8vSOerqyiyyqepZRSUlaVZdhVMvUvULKsqytRsvSrl06LHY9Cwp06KAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAgJyAyUpmqVQomamVZqlmWVJZzVLMpKiZZFCVSSqWUBCEKkIJFQIQoBKhAArABUQgJsAUEACoBAkEBKkFQChUgoEKAKQQhIlQhGvSeh5usc9UllVZRVVqUVVSUlU7LsdOyrK1l6lI9SrHY7Ksqx6FjDUeoUD0YUAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAQoUAZLNUpKonNUsyqVSysyks5syqVSoUsihSokSpEIQhCohCASIQCEqABIUCAQgRUKgABAISFAoKUFIUIVAoKBAIBCEIQhG3Sej5eufPV1RQ7LKKp2VVFpVjq7KsLKStStR2Vcuqsdjsq5ejoR6j0NQHTooAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAhCyAzVgpRZyUqlmVSqWZZlFnNnNSkqiVkUqhEiVCEiVCRAIQCRCEAlQAAhBYgFRCCkACAQCQURCFQKBUJClAKgIKUIBCEIVbanoefrnz1dUUllVVOqSqopKqrKsqx2OyrHqOyrHZVjsqx2VqOix2OjUKB09AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACFCgDNWCUlnJSqWZVKpYlSmbMs5qUzUQqlkIkUTdCJEISoSIBBCEKkAgEACAQCoEgIAEFACABAJEoigpAqRKCAQkFBSIQhCN+k7PP1nnurKKKS0q10yrKqikodlWVY6q5dlaj1Ksqx2OyrHZVho0dPUNQoHTooAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACJyAgzVkpoJymaWSmphLKrNJZzZlSmaiVmFKhCJUhCpCEIBCQAUAqQCEIAEAAIAEAqSFIFSAgCFQKCkKAQUhCAQCCEIRKJd9zr4dM+W7qirKKSiqodOyyqpHVJVlWOx1VjsrUdzVjsqx6jStSqLHY9DUKB6OgAAAAAAAAAAAAAAAAAAAAAAAAAAAAACFCgCDNWSmgnJSqWZVKpVEqpVKs2ZUpLIpZFKCiRKgEISJUIEkAFBSCEKkAgEAAAgEAqQAIVgIIVEIBAIQhBSAQoBBCClGRv0nZw6Rz3RVUlFJQyqY6oaXVFWOmlWVY7KsrUepVlXLqrHrNWOytBHqPUNAdOigAAAAAAAAAAAAAAAAAAAAAAAAAAAAAhQoAgzVkpoJyUqlmVSqVRKqVSzmqVKpVCWYFkIQhKhAIQhCEAgRQCAVIQCABAAgEAgEKgQgQVIAIBAKFSABCAQoKmIVJRv0zvw7Z8t1ZY6pKKShlUx1Q0uqqh2Vc1VWOyrmtHrNWVY7KsdzWo6djsehqFA9HQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAoIUEEqgyU0RMKVSzKpVAsypVCzZlUqUlUSsyoBRKoQSqxCEJQSISKAUAhCpBRCoABBBQIBCABUgQEAKgFAitUFiEoiVBEkwU0kiXfpno49c+WrqiirKGUlDKp1SUVVF07HZVzVOyrmtHc1qVY0rUdlWPUdOw1HYaA6dFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAQoUEEqyMlNBOSVZsypVKolVKSzKs2VFWQSswKoSiJUJUISIBCVAiEApABCAQCABBSgoAQAIBAIQAKgQQgEIBEkKoqlEIKIJtvOnLrny3S3ZRVjKKSih1Q6pKqiitSrKsqx2VZWo9ZpK1HZSPUqx6gVqFj1DQHTooAAAAAAAAAAAAAAAAAAAAAAAAAAAACFCggzVkpSVQoUsyqVSpVEqpSWZVklSkqhVMqgVSghCASpEqEJASoEQkFSOEIIKQCEAgCkAgVIKIhSgrCFQIBAKFbEIAqYQK0BCTbc05bz5btbsoqxllI6ooqqKsoqnZVy7Kp2VY7K1Hc1Y7Ksdj1KR6MeoWPUKKB6MKAAAAAAAAAAAAAAAAAAAAAAAAAAACELICDNWUykplKqFmpVKlUSqlJZlUqhKpSFUyqUFKlBQgqQEAhCEAhICBFAAghAKgQgVAhaghAKiAQgEFIISQoIBCUGIQEyTCrfeejn0nlt2UlVRRRRVMZVlFU0qnqNKsdjSrK1HY7Ksqx2OyrHqOx07HYaOwooHT0AAAAAAAAAAAAAAAAAAAAAAAAAAAhBCgCDNULNJVlKqFmpZlFUSqlJVLMKVKSqFUyqUFKKhQhUCEAoCaBAIBIgBCEAl4o4tXojI0Jrkr0cupAKUAlSACAQiREjgpQ6YlRJMIQDEm25tz3HLdJdjqiiihjpjLsodUjp2Vcuyh2OytR2OyrKsdjsdlWOx6CVqGjsKKB6OgAAAAAAAAAAAAAAAAAAAAAAAAAhCggCCVQZKUlWUqs1SyqhSpVClUqlmVKSqAkUqUhKKhQhCoAQoKQgEACASAGMutnFLuni6vt5mMu6eRp0BL3IgEoJARKzCEA7FK7ABEiFKgHSAkIRtvGvPpHLdJVlU1pLGUFUMqqRrVzVOx2NKsdjsqyqdj1KZdjqrHrNWOnTuSnoWGgOimFAAAAAAAAAAAAAAAAAAAAAAAAKCFAEEqggyUqUhSqJzqZVAsypVKhZqlQmiFCFaoUpCtAlQgFCpAIBCABCABAcOb26mEaoj53V+hzOM4tPYw511SVQgABDHYCVQhBSgpDABChUhSiIRrvOvPcct2lVVNKKKGOmMqqKspHTsaOyrHTuaHqVY7KuXY6dlWOx2OnY7DR0ahQOnQFAAAAAAAAAAAAAAAAAAAAAAAQoUAQQSqCFmpVBAqic1KpVKiZUpKpZgzZoaIUKlLKkKBRQQCiRAKgBAIQCAEF4cXr3GCTGNfMau8fSZkxVIIBVMFISoAAYhAIBQqBBCpQCWUFRr0xty3HLdWVTSiihjKoKKpjSrKDSkdjspCyrKsdOx6zSOx07KsqwsejR2GjosNAKdOgAAAAAAAAAAAAAAAAAAAAACFCgCCCVQQQpUqghBLMqlUqFKpZUlUqiZUDRCCJtUKUhKAqAUIQCpAAgEAgEI483s1AkYpPxj2Y+/83T6bEoQkShMAqBAqABAIQoBAKkEFKEIQhRr1m/LUc9UVVIylpGOmMZVUCUVYVVjsLLR2Oxj1mqdzVjR6VcunqNHTsdho6KLCgdOigAAAAAAAAAAAAAAAAAAACAUKAIIJVBClIUqgFKpZlISqEqWZSVSzKoUqCVEqpQSkJVAISiJUgIQUoKQAAgEI8/N9DWQYiY/JfVn7jhr6PnFSFKCpIKgEoAgRCUEYZbaAhAAhCCEIRt0x0cumfPVFU0pWUOygHVFDHZSOmjsdjsodjsaVo7HZVy0dOx2VT1kHqUGoU6KLCgdFMKAAAAAAAAAAAAAAAAAgEEKAIJSFBBKoUqhSqVSqEqhKoSpVKQpVLKqUiVUJVAoqhClVIBIgEIAFQAhgIBDRHnY16O8ghAfnvafXcr6kgTAIQlBAoiAQCAQS+dL6GokFBCEEgJQQjTpnp5bjnqqpGtFDsFoB1Q0Y7GjHTsdjR2UOx2NHT1GlWOx2NHpSPUdhTsdOwp0UWFA6KB0AAAAAAAAAAAAAAQghBAEEpCgySqCVQpVKpVClQpZVSpSVQglQlUpCqc1KoFFUIQlQIjzl0ILiKqutAQDQEJQAQPPxrv3kCgE/P8ArPpMa9vMQQhCAUAgUEAgAQHDNdtylEFQCRACpCFWu86ctxz3VMZQyh2MYDV0xyOmVY0B2VRZSOxo6djqrCyrHY0qx2Ox07HY7HRTsdFFhRQFMKYUAAAAAAAAAEAoBQBBApCgghSpVkClWaiWjJKoSypKoSqFKCBRSFCJUWYJUCqEIBGBjL1WZmcu+oDAkyhkm2oxgJPL579XpgpQUHwPV7WH0OBSUkBCgABAIAEAlDz8a7t5IKQQCAAEIC+knlvPlqih1Q0Y6cUMYx0DGUOmNHVWNHY7HZQ7HY0dPUdlWUjsdjsdPUaOnYU7CnRRYUBQOmAUAAAAQAAoBQAAQSkIIIMkqVQQKonNCZoFKhSypKClUIUoJQFIQhKoUoKVKCEIDnzfF1fTzOzUZIxERia2JdEqhA+QdPPzr7jfINhoj4To9KX6fEAEEKgBQECLsJQQ0QHnY336yUQgEJSFXmr8n0vzvSfL9Udcf0R8vpnz1RSModMcUMYx0DGMqmMaOyqY7ljsqwHcuqR6jp2VctHo0djsrQR0U7Gho6AosKAHRQMQwEAQAAoACAJSAUEAQRLQEKEEqlmUVQhSpUKUlQClISoBKQCUgEsilBSgCAD821r7zE7bJCiPOa45eY+T3fby808lfG1eCuHSxSlXHcnoSYdMehH33J6qdCddigFRBX5c6fHb19PJ7Ent5zR51vn15Gr6uZ7HO/Ta57Aky8h4GtfObfN7vy3R525NismvWuf6T+T1jnppQ6oYyoY6YDHTGUMCrGjoR07GlWMdglU7HY6dlXLR07HY6djsB0U0dhoUwCwooAKYAAggAAAAgCUCEKVQpVljnRGGN4Y3yc9iZyxmux1pSIlQlQolZGMuzSt7no1N7HRCUhAqglQCVAB8Rd+zzePNedb8+15i8lSiPP657uepWKmzzuk7sazRVFXE1KcfTOOp6HLaLjsl9iTvT0JPPt4V+a2xsRNFETUUIRNdUpL6Uz5W3DZNTSSaViEir1dZ/pf5PTPnqqZQxjGAx0DGUMCrGOwHY7GCVYx2OxjsdOxo9SkLHZQ7CnY7GFjp2FFA6AosKAAAAAABSzEyqVZTLGbhz3hz3xeftnLlnUEwiYmkqEiJJiCZUsErIiSISykxKzRE0KzWzs1n0emO/eeqzazo1NLFKHn415WN+TNeJnXx/Z081LnSIqLEqPM659DnqSSa4tzqzYrms3lCbJOHpnl3PU47kigmwh2oEQCoEiFarEgJZqSbEICaQgRVLM2+rvH9M/J6Rz06oYU4dAxjHTAaUjp0IWMaOmjoHY0Y7HY6LKR2NHTsaOinY0KY7HYUBRRTAKiMsbzxrPFzzrPGs8azxrLNjOolQCgCkIkUpSEKJEQqEiESRErMSskrJMSSTLIiRVKzCpCFCoUQGdOp0XOS+PnUWZWwnz/ed2GsTUKqmoFXk9J6nOwKoODpOvFRybnTmwRSTi6Ti6Z9bjuSAM6BWKiAQFE2NZsUTSpEWAhCtSIQURNiJr1tcv6Y+X1jGmOgaiVa0YwGCMdjpgjQpo6aMKEaFMdjp2MdjuWCJSxDLsdhQgXYi9R1z43yc+nPz3zct543GbQFI7BRJlVIAAQSoQhEqgJEJJWZUiESTCWSYlZJWYkRMSSJZESJZJpChVJIiQABCpEHhd89Wb0ZZ1JNk1JNeL2nr8bFImvM27spOLo6Odw3JW04dzg649nz9YsmpIpJKiFSTY4azYAJVYhVKFqQlVSgIKRIhJ625/S3zUY2DGOmOmA5HQNHTQriXzK7pM685eSs15TmtiMjkWI5VDGHHQkZtRUaRpLpGsXFVa2UmiOtI0sdXGiXV2UUBdUjSgBXVJZQDVgBJIlUIRIiVUkiJFCWRRKySswqmESKWREiiaSxSJiSaQoVSiUAYAeL1nTL05kGVKoqLEeJ2ns8bIrYs8nrPR52K4durFx1M6S8m8+X2x73m6SRU1AhUhE0rJAQrEAySbRETYKCQtQEoqgSepc/e8q+W4XdOyOa3QyOOzGuZeaucg41DmrzqyqjSWoouNJbkqW8tC4s0jWSzVN8t8t43io2l0jYsss0GgajqDoTGKTatKutLKLkQhEqgAcKgUto6YFDKWkqpEKJJEqFCJhEqiVRMIQpZJESIkki2SVQomxEiESMZR5PRvHdiTbBlqSZVFnh9nscqCsk8jrPR51nn7dmZnbjWNc+54vbH0fm6QTWdMikJYsiyomkAlmxE6jlYEoqkhZ1KhkVy2Fa5ce8+5Z5XXPlZ1cpLRUNXDHK0crAZcrihRctGkrLlqGXFwzSNI1jaNpN46MzaOerPB63sypPoeLrzeXSU9jF87ecjol0jQ6YouTay6F2s1NrAEFkiGAwEsqIoVIUqEAyhmllAIoYoVKEskqiYSoUIQiSSVmpiKlZEkiECSADUPL6NU9LnWImoIMtT5/vPZ42SSdTx+s9XnYPP6O3DOsKmubc8Dvj6Xy9JJqKRNSIky0okDg3JrtxfJ645N56s6CLOHeezOvN6Y5t568bzuWuGs52SjXHWfY3n0/P38aXK56sdJTWVLcsowAqGMrNocUtF5rKNM210y0jSKjaA0NY2k0jeTfL5j0XKiNo1jsjRNpN8zrwnTbLaXaXojSNZdE0soqqGaoK01qTKJNDUdBEACEISolSESImEsCGUlK7KGrAYDGSEIkkkRKySTbKTShBCpACJfL2VevzOHQIkivn+89jii3NJt8Xtn1eVk8zrO7Fyrm1Itw1n5/0Y+q8nTKvN6Tpzrh3nye2alaed0zFRZlWsuVkWMixCpEWAAmW5cEoTSQRUrPars49Ple/HDWN89EhKzpx02xvfGt86uLlEctQy5ai5aLluW0vNouNctI0i10k2ijOztw5NvA7KjSLjaN5Ok6My00jfM6Jds3aNo0a0NZNEqmUjLVgJKpLlGptVIxCAQlRIgWYRMoIgkkkAWBASIkkkKIVUIkYhhVwwJLAS1JNpIUjzNsK9jmZFKHbic2nNqetzcmnnbce55nVWXNp53WdGXldM9E1jY7PN7c+rl0z1ISaVZ6l5omeoAjlx1mlqWLmiKRNmeskTSscKosagDgI1n2tTo5b+Y6841lyg1CpQ1xr1/N6OznsGVLcOKlqqzaLil0i4uKjbKzWW00i05q8Pq9HleiOHo0hojeOvM6E0hybxvJrLvm7y6xcuhsaXNDLRq4ZJIwoLVm1miBIKkSolVCEKJUETE1JIomkqWE5Eit5aJJM6RNQSTWdCZrlqZKzDSQMligsCDPTm1N8XeOLSKQzeVRnUVz6mG2Gpz6zcuWs52BjuC1Jx9cbY1JRlqSkWIVgUpGdk2Usk3KpBYQrFVywlFzWmbpNTYjOzSXLU9fWOPry8aWLlq1IClReb1c9+hx69/LppLUXK1cWXDLi40lovK40jWLKTj08PrC2bNY2zdsrizSOnLtzNZNBVrGuZsu+b0Zmk1oVW0ao7GlRQNACQURW2aGlCXEioFCWQhVMIlQUJZJSaylgCjOuSwl6Ea4WYUhLNJHHPqxUmNYl1Bw6SvRJhq41FaRhTCubU7OeosKzMNJKjaN82KmxGGnPqZ6ZXOOpnZFKx2cm81LNOIsAI1IRnTnUlxrNaRjZzbwqcuksHRnW+dVlnqC8u8XAvB25cfblpm742j0O3HLWPFlAGrla3mqnDHL7Hm7+x5+1ysZcUOGb5qNI2zdZNI0HHn7nbl8/2nD1zebtLrGkXLcbRrHTmbSdEu0iNo1Nst83eNJbqzWNUpKRrcJUKnE1QAb0gjSxiGSChJMZRlKq6NTY4s6yGSYgSMZz2RVSqzFc7GWuaZaqibM7SOfTKrgPO2VKObVZFaRFSRZlp1YuWpBhq82stYSjfNtbyiybc7Js595zNFRtCPO7Y6uesNZ1zrSXg6Yw1l1NjEkG2d+nx6ed255azvjXH15laY1hvAIqWNSSdZRNk0IrIsD27MdY8aUGoOVl50AOWo6+e/oPL6OvG3FijSLHLRxab4dmbvmdUmpznynry8sttc3WLi41luNctY3NJN5N5enM0yK0OjN1y1jVaNDWNEtGNagJpFCJHQaABYhRrWZMJYJJhVmu1mcsERVOoyKyM0pZslaRrAjKoMaCKxshcqyqBW8O5y6XARbUlSzXNpnppJGhmxqIz0ySybLWUua0y6c3pxZrg3mbOrOt5Jl8bvjqzrze3Pp5687plkWYdM741cqs87txixBV5sWUtSuVWZaxluARcs2TYKyUKcRqOA9xObrz8WUVgripalqUHFLpm9/Lp9V4vRydI8uXedZe/npylctb5etydmXRmM+T9U8vrmpbluNI1i5dI0i5N5d5N8rTWN5bk2XXLeNI0l0LLNYtLgGNWSFgAixUCGrhgXZEQpYpQYoyMrZEIIRIGdk2sQFmJho4zszMNHKjk0zoXI1Ma5Kz3IMdOzFIx0uMdLjOsNMLLFSosUSYamkaqjM7eerMjPU6sWLGuOmes+X2xWLzbzFcnXmrOrn0y1nHWVcpahVFgRqI1xoRVNk2Kpsmy80WNRIqBWShXvRlrHiStXKylIqWpq8gCo7OfT3PN38X0cUTZpLcvocenqcdqXoy9LDTLsk87b5r05iqNM3WNIvLSXQqNo3jeTTMs0N5dY2jfLeGukWUukaSaIwGNQQUQqCh2SECsBGgyrBSClGEYGaySTY5QkInUmplVaRcuGpgKubUzrCujNwMNJrCmXGdRbknH0RWmXTm40iNSBy46mOmWoFS7xK4aykVudOSK1lcqibGCtKijm6Tnsz1ETZz9Mox3nO5uWpBQcs2Z7zJGpGsuJqNQFYRcumdZazNisQrEhXvy53PiDmmOVq4qWoqaBxUuuLrNTYFRS1L0Y318t9nPW+NdMm2WjPzvpzNumTNJdIuNs2k0l0zdU6crk2hlpqvTmbxtLrLtkyy1qNUuGEOgQAAE0VY4mnDGSOqjUBkGZjLjEaTCpQqZBJJjpmhays2LM7IUSTO1pz25VjphWkOOTogqax1JpyRWdRUUi4mstCEc+81K1EJSzMaOI1MxkWlk1ti650iNZ5+mXCl595Vk0kmpsz1nLWVZGoLUVKEakWOJqxJU1NmWszYxyzci56xTXuxnceKooMqacVLebpnTRrJpGmdKqhxU1a9HPW2Nb5vVjVx24vm9ccfTNRpLpm2txcaRebZ0ZaL0ZlFSNNTeXok3zdpdY1i4souXQuQAYxKh2AhUURpEhVZXUgMmW7NTnljSYwyyqKUjtCKuAxrOsqys0lYozsikZ0lxpGdYVlUVlWeihE1JFKpM6y1ENXJFXLhrOW5JlqCBpnV5s2Z2KzHUcZ6m2dTSXTLaXbNCs1GVnn9+WO5Gs7Y1Fc/TnluMSRqRZct50yLEmudVKrCVWc/TnNXNXm47xU0JpnXuWcvTl4quUFY5Wuma5al0yvOtc6x1i5aWoZ18ums1eVTVydfPXZnXRmfP+nnnVGudXGuVq40jfGtC5NZdpNIcXZpGxvJ1Yuq6xpFxpFLZcXIKqpGqgpWVLIak0o0HCDK9OkyrnhS2mxzLkSYmemdlS1GdI1gEZ6YVFSZWJakRjbzamdqJqTK3n1IMdwBbyDj6TKs9QhLNjKlzuRWZaiSKFyuZ1JN8aqUskiwMtSK2zal1zejGsNZQxCKEuG846zjvOHTnGplqMqWbEm+NTUWBOpeNMqXfG+bpzmwViSdBIs91effHxKctSpSqlqW82oqWpejnubHGkrWLN8a6MbuVwrPQ49O3nebpnyu/PTNZpLpnWkM2ya9GLrGkM3yLLjaGWnZlvG0umWkaRZa3lotQrKKGshUI5SxCISraHFQ6uwjnVRJZz1UZaZEUCJMzWHUGQ6Z1ZvLqYaB2ZedpzWcm6ltNIzqV5dObUy0uAcZnH1mOpJNKyRxUqoJuUKpKlI5+mc7GsazWaQquXbOps1xYq5YuZqRjlvN0W8sNTHpM7nn6Y5+vOLCpKhWVNOGZayqcAFLKTokuWUy3lkWe5Yk8WUGqHLpKRpnSqo0zqo1xrSXXGiydOjluyAsVa41pJlqMuXSW5al0iio1l1jXN0yo1h1cmsaRrJrG0dMXLrm0lLpG0XKwGUMVTE2CqSKBIBSjbNK0rMzAyAVZpBGrmjWDOqiUdVGVsaaZaxNBhVHHuTLuZmNdOb0ZY25WeV1SceoxVzac+5nZIVFkahlS3KyGRVU04IjUw1nHeY1HmlmmdaZ1pmhNiUEJMtwNM0Nc6rNaEsaY7wGepz9OeW8qhERqOWbkVWTYwFYhBUoybA9u5JfEBWOVy3NJGVLUt5tS9fPemK5VYFy7ZtSxQbZRRY4Vty65rWouW0qXWNM3SLiltKjSNY3jbM6UuXow1jSVlG0bSkA6cjWNJQJAVQyKhCNJbNYyrMmyLUBmmVmNCpc7C1RjqbYdmb0wqztRB5+4zqzQwqQXzekxp1yaIQSYaAGOnL0mdk2Vm2uWsouWpcrI1lSzZNOETZGpNBti5ammakFSxc57yLFkWKwLzWtS3nSBGtRebGplrOPTM3OepGsxYLnrFLNiJuamlZNjlVyKCRnuJFeKpDVysauWs2hy9XLprmxc3nWes7Zrloqa1xaUA0ipQdKrzbloI1lZpGubpK4pKl1NJKOnM7+boi4vN0RxpbUaS3FDlVlQkjTKmMQibCEMiqNZWSkLFkLGlyTEVlZnq5rFkLFKNZPQw9DNDOs9IM7FKyK1luCOfblOfTn22xbIRrtltGep4PeeX2ztm65uNmOnVm+ny14/Web1xhvM1CRqOBVYpKW81iETU2RrM1nrKAx3lrUIcqscpQjlvN0zpysmwXHeMt4myNSbJsVk2IVggqQCgSB7tTHiytXKWVNVKS1DLzejn0VzKCtGoaZrW82pWaZt50WbZumdaSqwpF5ty3FW6RpLUCXFmknRi9eWmWyI6cqzas2jWWo0lDSCqkmsKz0clqhE2IUhQomjVRKBBnSqpYQrOsNMKlc7JlK0j0ObckmgpHBUVFkmN1nZkudZ1nWdTWVZ1FkjiKmuzF9Hlri3JPY5Pb8++Pb4b245OmOPpnPWctRCsFJOnG0OWLAjUi5ms9Zz1lW1E2RVyhNk2OVgIcdnLo5Zs357z1IrHpzz1M95lI1mNZViBBQBIrAViPcuXnfjzQpANXCs0zqpdsa0xrDphwqqBaCNJXLebS1F51pGudCU1ti6zTkw3m5q40lqXWHQXFxrl14OXVLizpyqNDTLfKy4ChrUkVz6lgEO1JBIkAtK0ipbkFySKVsWVLKRXLphpnE6pE1vl25aJNTTjGubSLahjTSWkztyrCsajRQqmosmpMqzrO5RNBeb1ZrzZXrw8vvnpylNprl1nh6Zw1HLz7xpnU0kw3mNZVRZNiscrIoRrFhSQActRedBRvy6a5uWpj0xGpnrKJ1M9YmpuUgIKBWAkK9tnbn28aaCpRJqocpV4ty1LlrM6lZrWoVlZ1RebUty1FS3KDW41xqjozqouGtxa3FxnqXFS6R0YrGmkukm0txZvJ281RrLKLSoqIqLLhEWyKylzEjS5Zt1NMgzsw1M7ZWAEirG3n0zETVr73F24vbHPZx7nHoji059XeOastBNI1gMLefcxsztYrERUgSZ2Z2RqZ2CouLmtTk1kl9Dnv6zyb+g4a8Hd8Xvjy+ufI9HLOyLMd5z1JsVkUE2VK4jUByxrKoBHKqqKlFm5DXG9M2amo1mblLGsZ6iuUKxIqASbAVnumvPp4q1nTUk1zpCsuavNz1I1lI1qVAVDVxctZumdWaY0qoDTOtc2zXOtsHFK6cs3O2dCXK61y2zenKLNIuXaGa5dmV5dWVnPqKunCakysk2liqM6RcJLhWpFTiKxrLTK2BCGRWdsVhYFG8byXL05txnpz1nXLpcSc+gitSWtRrHHuZVnpIrIHUChVFiSNM7IslZsAl3jt57495w1nTOvv/AJ3o9Xk5a/N/pcODriNTLWct4mpsmmqRq5FUahCsFARyzY1vIVWRqEFOXTOgDO5nUmwSNRIrEKxXKAVnuVpz34i3mzTN+fS86z1hrUqJsLEjEtQ5QC5dcaqVppndLUM3xqopal2xQEFE0XozaN869DD2OTTN6U8XVx0SaS6SUejzKLiaiqNspsyCorpyYCMdFDLkm1VFjHm46c2mdudk1KuFU1CZ0FFgWA4RFJaIrOxRSpAjTSGY1jUkakhUpNKFU2STZFZ2IjUhC1Cro53pxv6Dzb+Y9fLu5dPV46+c9GOfpjDWct5iydZz1AmnDUQXPWWICoFARyqxE2KlYkVA5po5pJOsuBZsm5ViFcqkir3UedeLLUtTaubzq83SalGqsQI1QAXKhJ043Ixx9L5O/i98IuXTNZpLUrTfGosa9OX0HHW0XL5HRvhnXs8r7HNnXJUVJx1onfz1nZeU2Z6bZUkrz6RVydGW0c9ZaZVnbcUaQ0KRkXHPq8u0rJFgjUsChUCM9RDJJXTK1ZzalwxSuqknRxFZVjYqipACRWRSSamyKhJpEak2SImxr7Pm6Z0LjqVz1z9MuMdTDeMOmI1IsVOWLmlcTqSlK5QEQ1mybAViSbAVIapkGtTQOVWJJsVyrJFYrPdZed+KOa0zoBahyuJ0qLzpIqqBZs0lIpfZ8no8r08CKl+h8vbx+2Vc1LtjSrozpxKUqTsxr3+GiXj6Z6sXm1ePpHm9mHoc7ybntcktdknjbkr1YdMEc2k2ONox1dZA1jM65PP3cdMazoLlpNYRtGFm8ZW8mmVTQBaWOFYrZoQM6ioGVLUQtFwGg0zqTKsrJqKiyFEVBNIVmdiERYqkzsnUkCbIsBHuebt9N5O3yPs4hvjUy5WeZ6OPP0xGoidQI1El5s2FVK4FBIqViRVNiFYkKIBWAhq4agArIuUzNTrPuJeNeJakctTTAJblEuaSOaaOVgs3OmdaZ1rjUazUtRtjZQm2NVK6eaWA1cejy3rHJuCTVLUu2bRtm65dOaR3ZSmVQa51rJnVoQwoX0+V1Ti1OXbOuTaQW0lUaQJ15Z1cUZVlpz6lRRYRoSdEcuiqSKRUVm47kW3CTSGsBZmY7mYE1FkqGdisQSrUzsCUVZ1NlRlpNSkWCKkTZcv3vzPWTV6z8Z7OKNMaw1Js4+3Pn6c41JsvOo1lWOLzoCxAKiFYLNkawSlJJuRSxAAIKwHK1JVchNis9xHnXiDUAVhDVxc0FSqwlvNa6Z1rmscEUvby3zalyzci743nqXm3K0BVUbZ0yyUirl0l2zblCoZ14vXjXbmctcG5tLUBtkzbLcZUUnRl4Pe2cupFawkGoCzTLojGlXTi+nzTXNucmhZR1YbS8umFAAWSYVjoxFFxRmRYLlZz7zNtRlqSIikTYwjPUmxkVNkUoVRZNSk2ICaVhHVjf6J8r1/Q+bf5f9Xh5vbk5ru56WNed6OXJ25zZjvEaiQRGmdKxIKqBWJHKVnrLlVk3KFYAiCiCgSNXK5QLEB7qI8SULlmpuQauVy3K5Z1kl1xrp59M9ZqXTNcALpm751jqUmdXFS3ndRUrsiyhF5tFSqmbZuma5dZXVRcb5vXi6ScejjDS4uKN83pyaXG0udeT2y1SZ6AErFVG2WpmXXdzukduXl9J1w7Lzbjn05qwqKs5NzTNy1NM0sI2WoyqKknSY5tRWUI59RWZ04BUrFLlrKqoz1FSiNSRGdiqblDJJsBV6vn7fWeD0/Mezh5Hp41Hbw7d3Hp5no5c3TG2dZ6mG8Y9MRc6ZqRUgpCSdRDASKkisCbGTYgGJGqQolauFY5Q91EePnUWMqaz1hJc1Us2VKhUzXG7zq81gBebrnWmaGepUojNM9KhwLGs3E0GktZMKuW83XNa1Lvmqkmsu0dOLpHFq46yAmmbrLtmyz0y9vNxdHHtGmuZhoWC0Z10870StM6Dpys68XZFGWgZHFtpGdcXSa5YaahAtZmw5ZqKysy1IM6oRnZnU6kxNACJsmyLBSs7m5rO5kiwqKlFZFgqsImxVJpNaY16HLp189eR35dvLplqXJjq828c/XE3NwhkpnqKlYQqViSpqbAmybksBCRWCiCsSFIYoauVWe4JPGlByqlc3nU0I1cADmmVLUrlcty3lcumdjIqpwFSs0zpE3Okuk1KJWVAazThmmbpLUs2bS1FJ0Y1mu5yamVjLluHFHVi92LvHB0c9mWmdkajWzSKlvKjSOzKzok2xrl1OTTPSomgxrl1CtcqJrXLaLjKsNGYaIzrGygMrJpEWRYwlVTcxU0kFixWEok0kms9ZmpRE2NZsSKiWbOrG/ufl+z0uO/g/p+XbOsemPc8vbz955emfP7c3GkvL0xNVHP0whWAkVBc1ncqxWRcliBEFIYkFAFY5VYxDl9rWXl400rBXKI5QVMIVjHNNazalALzq5byqVgok1ea11xqNQGjluUSpVQXK5ds6uGXKi41lDWNc0XTLj3MtRlS3AaSdWN6RtGVuVmGxcuHSoGBcukehyvr8rwdDhJxbVHNtnXPqNNMXaEtlG+WdQZalRlq2nHqZaCBnWdk2Cwis1lgVZayRNNYsQrJqokiwrO5mkiqUKlFU2OWLNJfR8/b7n5nt+Q+l4+Pc9Ph19Pz9cdZ4uuOLpnn3ibayx3jDpiLFYqFIm5VTYwXPXMASFSMVySrUJVY4AVWA5Q9rWf/8QANBAAAgIBAwIDBgUEAwEBAAAAAAECEQMQEiEEMQUTIAYUIjAzQRUyNDVwFiQlQCNQYEIH/9oACAEBAAEFAsv1f4xXbL9X+MV2y/V1X8XLtl+r/GK7Zfq/xiu2X6voX/rb/wDALtl+r/GKMv1f4xXbL9X+MV2y/V/jFdsv1f4xXbL9X/Vv+G2xXWX6v8Wtl2bdF2zfW/iavTZyzbo2csSdZvrf+0r/ALWyiq0splVou2b638TWclaWclelds31qKKKKKKKKKKKKK/hazlm0tLSjb6rOWJcZfq/wXPrMON4fEH1cdvVMyLqYLy+pP7qBDxWLz4+qw5fnWcnBZybfVZZRWqMv1v4IhkU2dXCM8MMUca6mD6HNCSyR6ith1/VSxHR9JHo8PV4oTj8izcXpRRtK9Fos5KNq9aMv1f4IwfnMyco6Rf4XnOr6mHSYOg6SUCjLGU1yWbjcWzkpmw2orSyyyzk5KNvzcv1f4Iwc5PRlwwz4peKYvBzo1+J5qRts2opFa0UUUUbSiv9TL9X+CMP1NO+v/6EezjvwP8A6FGX6v8A6y/kWX6b+ZenSt+Zfp9v+nnPpvAMM+m8I/05Zowl81GX6v8ABGH63p9uF/g/DXu6D/Tzx/5vnZfq/Ov/ANR7/ga96xk+txY17zEl1cYkeoUsnyK1ow/U0rX23X+C8Fd+E/6ef6nporWvTl+r8yy9bLL0svWy/Xf/AJby1thPYNWpyWNY4uQ/Q5KIsykb2ebFNOyvRghslXp9tl/gfZ934L8qta9XU/U+TWlFaZfq/wDt5xo8R8TxeD4YLzda0o2/FOLxttJY4MitK0n7T9LCcfaLpty6jFJe8Yi09fbRf4D2a58CK+TKcYEZRn66Op/OlxRRRRWr4XUeJdL0pk9sukjHqPbXNI6z2g67rCPU5XHL9X/19fJ9tcUvw3pItdPRWjM3iHT4IvxrolCXtD0cTp/aTH+Lz9qcCWT2slWf2m6vIs3i/WTF1mbCtr0ssjmnFw8U6qEum9oet6c8c9ocvX+GeC+00ej8Ixe0fQ5IfiXSD6rDGeta+I+0PV9P1fW+I5+vl4D410/h3SdL7XYZv+ougJ+0PQQWb2q6KMZe2GDZ/V3VV0PtYpH430mZ4skcuLR8E+swY1m9pvD8J1PtrjRn9r+tymbxDqeoHo9Ifky/Vr1V8mvTX/c7kbkeZEn1EIHvGI99xEvEYIfiUj8SkPxKZHxHInLxORDxOo/ikT8VifiqPxZH4sj8WR+LxPxdH4wj8YifjEBeL4heK4BeIdOyPU4plr5NaV6Pa/jwafi/TYMT9pcdZPafKZ/GOqzqXU5ZLWP6161xhbeUcqOTdelFHXfpfD/0uiySi4+I9TjMftJ1+JY/a3rIkfbKe2Xtb1jMntL1s55s0809zLL0vXcy9I9XmjD3rMyfjvXzWXreozj1a9UPyZPq6UUV/wB7ZvR5kTzoHnwPeMY+rxj66JLr2PqMjPOmOTf+pZfov0W0LqMqIeJ54EPG2Q8XwyF4j07F1mGQpxl6M3XYMCl4708TL7QyMni/VTfjmfJk6TFzhaK5aKK1j+vaKKGjF9aihyqdaVp1q/tfDv0tfJv5Nav5kPyZF/yUUV66/wCuc0h9RjQ+rxnvsT30fWSH1eQfUZDzpm9l/wDWWWWbiPV5YEfFeogZfE+oyD5GihxPGV/Z4FfT0UbbNptNptF+47eKKGjF9eiiUf7ih6UdZ+l8M/TaUUMr5z1r0sooooogvgyfU/6SxzSe+KbzQiRywmb4m+J5kTzInmRNyFki3uRZLqccCXX40PxBsfVZZHmTevb/ALW/XRtNp4xH+y6WP9q4m0aNptKGiv8AJ1pRtMS/udpRL9S0OO0S3lHW/pfCv01DXprWtX66KKGVo0V6K1h+TJ9T/Q6nren6NYvaDw/NP8T6RTl4z0MTJ7TeHY5y9rugjl/rLoRe2vTVH22gP21P60ys/q/rN39V9a2vaLrtz8f66UX4t1ciHiXVQPxLqR9Vmm/PyM3yNzZd6Isv0XombnpZZfpUmjezzJHnSPPke8M94PeEefE82J5kTei/+ior5/iy/sujX9rtHEooY0dxr/K7eNtmwcaMX6uiifPU7TJH4McKxJM6pf2nhCvBtNptNpt52lasoooooZRWtH29NFFa0Qj8HU+3E+l63+vsIvb6HmQ9vsG/+u+i2/170+/+vem3S9vsNL2+ltj7e5kZvbnq8kJ+2viEll9sPEsh/V3idL2j8RUpe0PiEiXjPXSJ555mKTRvYnotF6UxCaLQmJiEfaE4yLSNyXrUk2JpjypEHalP4vMsjPjzDzBSsT+aptHmyPOkeezzzz0edEUk/n1/t+Kfouh/R0bRxNptHE20ZF/ldpQ1pj/XUzaZf1NGSHwYo7sM4vzOsh/beDq8W0rkqytKKHxpWlFejsL1OUTvo9MmeMDHmUyXCWdNwyR2eMfuyiUUUUUVpWlengrSy9LLLNwmznTkrRURItFoTM/UeUZOorpseVweXqnOUeoOl6jzSWaKXvdqHUNShkUo5su6akzzGRk9IT0Qi9IM3CZfov5+5nmyPOZ5550TzYnmRNy/3KKK9Hif6Lw7notKKNpsHAyx/wArRWj7Y1XiBVGX9VXM4/BhX/DNf8nWcdN4LzFxKKso2lDRRSI9i0KmZc3lmHNuGPr0T6x7sXV/D77FmXrUlHq52uuidRm8yUZbZLq5RlPq5zPe8lLqJwcsjmRm4nmyZZj/ACeL/u0sige8JEZKS8xFpHmRLNxuN5uZbLLE/RRRRXOiFonqkJISEkIR1GRvJvbWiZiySgXbiIWT4EIQhaIXpsTNxuNxfLfO4Uv9Xc0eZI86R7wz3g94R7xE8+B5sTei16aH6qK+V4n+i8Lf9l6KKGjMv8ptGiiiH7iMz/qtxOaSwTXkSzRcutnfTeCOjehzgj3/ABnvGJmbroY1+JyteJGTxJk+sy5H7xkS94yNKckR6jJFSm5nY3PV69yiizucHBuRuN43pj/J4z+7Zm9wp7XKbk/MbIzpvqCPUHmql8RRRRRtK9FFCEVqkihUUhHA2oR6fqI5Hjyb5dbKWNye+REWkSuUXohCFotF6kXpZY/9V/Ns3s82R580e8zPepHvcke+nvg+tR73A96xnvOMXUQZ50Dcmb0WX6PEl/ZeFfok9POge8Qp5oRJ9ZjhGPiMJPLLd4jOW0y5FGL6yG1+IRcMXWR96l4mT8Tez3udvxKVTzTm8fVTxwnmke85MqwTeM3t6dy+LOCzgiWI3jkLJZbGNm4sutLo3m7S/TZuLMb+DxWf+Xm90vWmYJbo0Ucm02m0ooooooSKrRCRtFES5USE4zOpzQhHedP1DU+p6j3iW3Y9tlKlEjAhjEtKI6IQhaIXz1/pdi9Hzqxs5RGVr0XpZxo0fZxPyja0ckWkbqXmUeczz5j6vKe+5kS67JefrcuXHh6qWPEuryMXWZIjyTb3seaV+a2Q4bclOUm5MY0ONlUzuJcuyTN1EPzREI7DPu+HZZd6dh9zsr9CWnc5JxRtNjpYiOBte5yZ7u6jgsyYdhHBuU4LGQhHZ4y/81NVL5GLJsF1KIPetvNaVpRRtKNokbTaKJtFpxBZuouGPJtc572kIiJ6ITIxLOBrSOiELVCF81Fm751aUUUPWifbRaSlQ5m4b1oc9o5m6l5w8m5yfG5knymNLa+BzLsx8mX4ZKG5ZIpKIoqlwk0xtRN6ZwJ0b92m6jcVY0SKGtWkPgh+ZcD7dzuNaUNHGkcUpnkStdLJi6GTH4ez3WNZUsZjcJymo72rhGMYn/FE8yB5ka82I+oSH1EVL3w993LK3Ipo8xyF1DJ5FIxv4PG/3n1V6EdJMrSjaUUUJWKJuSI8iXG0SKFEfVVmyqE45pUtFohaIiRPuJWhCEIXoQvlI7iYiyJfyWyyzHF5G8RJ7Zb+d5u9G43ElTLLH3aEtGOVEXZJKRtobR5SNiPs820yS3Paqc6N9DkqU9OGbh8qJdj4Sk0TlZY5G4UiORnI7HuHa08scHagKCR5J7tw8SMCjKUowUtqUtsS4RMs0fmNnwQjteWduHUOCllbIdQ7fVRcZdR8UmspJb4U8ajKW7zKbyWbzzePNN452XTfPqoxr4PG/wB5+XjMOVSjpRZTKei+IymFUWRVqMKNhmzeRHNleXJL8okLRCQhCKEhKxRsjUTh6JCQhaoXzaOxYiyxG4ss3G4svWOR41vY2WJ6Xo2PR6UbS0cG4kzzGiU7LLScstDk2WyVn2yctiyEtL0ldXevYsuRdDmN3psZ9tIyTNsDZFHlQJ5Nr94IYvMPdSfSfDKOWEkrj00d2TqMM440rPM2ucjhST3CcUTyok9HpY+TstxwOhli7FD4Gyyyy9L0sgvg8b/efSta1TOmdZIqyedY5e8x2vrVCUetQs8JJsj3z/nivhx4SkSWnUZFldWIrRIorVISZFclERC0itF6EL5163p29NFG0a+RZdl+hM4JsZuLN5uO6fCkMlwbnoz/AOpLmfCUqFFOMse1bqNzmpR5XKdKL/KJknYkeWzZo7IrjhK1cZbZb1IhKMDL5TahA98yRPfZnvUh5WRy7skfhnKc23bcu0rERok+d2telabjcOizebzdfosu9b0x/T8b/efmYXy+r2Qnlc3el2bjp+ocDF1NvI/iXBHLQstnJl6qMTJK3otEJ+hCIi0XGkREX6kL/SsbsTsqta1bobH6L9FDZZYqkOiydJfZrS+ftJnYsm7IqiyxpScokkUQHksbQpEpc3RJ8Wxo5Wm6iGbaTlubZY9KKZLshyo80UixS4XDj8WTbTbO6WMcTbzyMSFE4L0paVpu4TOw36YrVr1Y/p+N/vPye2qY9VrjE6GQdLzDFPnqcnl45TLtLRaIQhHYiIQmiyxERCE/Sheqy/RZYtb0rRF8ljejkS0fossZY2MujebqGzcSnwpFjXG04GrHaHpF8yZKVikORem4sslKjcbxT4leiZIsUzfcbOxuHKiLLPMPMHJaN0bxM3m/ncSTIwJDsfBuFTKHwM3UbzcbzebkNx0fJw00KKrbG6R2Gy+bs2lD1x/T8b/eflKN6L0oqiHGkXZHhQIx2HU5fNlrEQtIvkRdi4ELvohEXxEQvk38pPR6Jjlp9tw5EXek3RZIZdl0KWjLLGNaS7FG8vmXJ2LN5Jjdm8lIkxy5cje6crEMRuN5vNxKQ9bNw9o2fYujcb2eYdzdRen3ZYp2NUbhTFchRZupp25DXEk7aOSPZkn6H3oid3WqK1ZQkbSmNFCQiD+Dxv8AedH6Fz6Yw3elGKKZsKRRijcoqzYoyfCyS3OyxaLnSOkT7rRG4RYu6EIQhehC9C9N6PWx6oW1n2slKyMhSsySsixsvi+WyI2ORHkqizcUOOl0ORvNxfOX4XvHPndwnzJi5GXxYyxDJDZY2XpZfF0WWMbL0oeidCaGWMfarEd1ssUPiUnjbyNvdRuNzPskeTY4lEih+juUfb7+hC7vaOJVDIuj77tYP4PG/wB5+QtYToa5ohHe5raIhLn7wLIujHOlCpLNl2rWhFCQ0dhO1tIpHIuxtZVFikJoi9EIsTE/lWWWWWXpZvossh3m60ZZuGyD5k+bG9LJSGyMqHIbNxvsi+dkamSiyEIjhj2ufOYWlfF5R5cqWNkoMcRRKO77EmiRZelj0slwLs+DvrRVqtGyzcWWLSueEWWN6M3COyRY0bLc48yjRtNpRRQlpuO/ossTGXouCTLG9Mf0/G/3krSihK/Qj4S0J3pDs4bl5dEIndti0jI81xHJsWlkZcJlikIviMqN9lidssUjfxonzFiYpClqmWJl+i/RZZZZZZZYmWLhSkWORZuGKQ527NxuNxejlzv5s7FnIuRqk83Cy0NzeOD2vJl3OOTDFJ4mOcYzx5cbIeTkfuf/ACZscMa+Elj2JsTLJ/J2iH6LL0fooRFa2Wbixy43G4TZuNw2bhOh92rahw4UND9F6d38hl+jH+Txx/5m/RZell6IqiMRnYuzdRuFKi7GKOjK07CFqtKFotE9KFwLk40QrYuBCR90L0XpZZuLLL0sssss3aKdRsss3Fllkmbiy+OxvNxZAXIhtU9khY4X5cZE8Ut0cUr8mVzxUvd3OXuUxYXBS+GTXOW63MbcnY5OlwK0JNvJBx9CNptspop29LGWWWORY+RiiSxJRiitLLG9LGxyLLNxZuNxvN5uEyy+WrGih6VY9bL0vS9L9OP6fjf7z8qCGkbqN5ZellnfTcWdi9GjbRet86LTdpfKIikj7wRBaKr+9jnQnpuLLssssskyzcWWWWWXpZYmNlljZfobGMss3FiZusw8iiUUUOCHBI+3mTR5sj3mcVHr8sVLxCVvq4MjkxbJPAY1iU2umi5e6tSx9Nuj0vTNrosMpQwY8Jk6fBIn0fweS7h4fmzEvD8+PFDp/h2UYcTzHue6OXHsJaWWMsvSyPqssbLLGMsvS+LN5ZZuNxeljKJIZRIr52P6fjf7z6b0vSrIcG4vVuhSLEzcbj72WWIRwUVoiy9LvTdypCE9IxEyMxyaIyd7hS4siyy9bossbolIssvWy+bNxZYmX6Hp9i+ZFjYnpZuIMhlpeYjzePPkeezzzzzzkPIm+44jUkPcOckOdjmWh0bUbSmh2b5RfnTPPk1vacfEM2NLxSUo++Rlmx9VGMukz4G8bwuPWdJCUc2Ly5ZOmlCDGP0dyi9LLGy9GXq9F29NnbTC1c52I7nIx6P5+P6fjf7zRXyIutH3TGy/Ui9LEbjdYmKRuOHohaWJ6N6LSHKsRZGQpDnucXSTLEORZuLLJSsvWyy9NxuLLvSxPSxssbNxuGxsYyyy9IqyC3JtV2QlZKJN0PkUnFObbWVnmG+zuO9HzpZvLL9DHpbN7RvI55QPeckjz9yXWYccHGOZrBjZPo4Ih4VKUfw3I3k6ScH5LRtGR1elj+U/VZuFOjzKJND9FFfMx/T8aX+ZrStK0ooihl0X6b1Wq0vi/TEaEihLiufv9haI37SI5MXOm4sTciD2ndIjHcSjs0WvFncfGnch+YaK49DG6TlY5G4cjebjdabN2l6KO59GlWDCmPpIIy4eZ4KG6GyaTPyGHJCCyTjKd0bhTLFIlxo2NiZZZel6M+79EcrRGaJ4v+NwcSMqMXUrd0fjeLHDpvEum6iMovq8vVdH7tLKuJ8sbH8pDH61oyxSLRxq/RXysb/4/G3/AJmyJYmL4jsWLk7fM+4jv6I6VQi+EyzebhPnfZdC5G+YpykotmOEpuK+LTmlwoSqeSNuEtpDkeZ1Kdxg7lKQ2WSYtL1+90Wbdse4kbjcSmORY2OQ2bzcbyxsssRFCltF1M0R8Qy4heJ5SXWymPNC/edxudqTHk5vjRPkTodIY+G9Pv2LGyxiO41p2L1txJdTKZ02DH1E54NjuowyVLH1OKZKHTdas2HDjfV/U+zL0el/I+3o7er7XRZZ3b5WtfKx/T8bf+Z0ei5Hp9tX3+RE+8WJ6o7FjZYtEdtEQxuROG2cYSUsWHHm6jyfJeCGWD6XC8/UZsOwcXHRMp3Hhvgjy7dylbojwWbxyNxvog+C6bkbjeWWOXCm9FKyuHGyyyzcbjeWWXqtG+Y5NsfNsi0N2Vyki0m5Wfdlj7VS5I/EfZj9F3pXLL9L1vW6IdROJDL5g+iWLBKTtdV8Gfq455ZPiGMfqYjt6O2i1a+RZZZZY/mY/p+N/vItVp30vj1fetEPHSQ2I8N8P97jNbZdzH3oTO5t5TJS3aPldNi87J1nQqC6TD58cOKPSwyvc4ZMSgsrUen6ifR583U5c50rxuPWdPMlgxSxdT0nkCE/ijKn2i38V8bubVdhyUxqURz0jIviUhz2rfS8znzDzBSNxuOb3m+1Mssb1vTbx21fobFIjI5P/nSxuyK3a3RubJPVl+ii9L51v1qTi8PiObDDycmWC6TJPGt2NN2bWxYHUsfMoUMetnYsv/Z+z9eP6fjf7zonrYmWP0/YZ3OxHiW7fCXDOz8O6tdFF8kStKEm1ZZfFmPJLG/CnGPV9X1SllxdTIXiG4nnjki8jYmTzWodQ8UcTbH1kpdNjn8C6nz8s2o5XPmGThPlTJSEXcr4T2mKblPJj25fJTIiltJSJyNxZZuFIchS5crVmN2slslSZYvRIrna9K0b1pi4E3FWJCF2SFwN82b7G0Se5svTvo3Wt3p3OyEdvR9itNx0HUSlPxiE4FZFGOd5Xn/t8nnqTyEh6dzsWP0ff/Ussv5GP6fjf7zrel+i7L9C0fdFWLs+XtIq9Gff8ruy6FLhM+96Yo7ovKqcjdS3cbltsgMclWPLsbyKT3bF0/UeWZMnmOcHjccp5gp0OVn2TLKMNwyZ445zUdksvwNZeZTtWOWiVrdRY2R5OxIg1EtRMqteW9rjQon37Jcqa4iqbobjclT2EkeWRxNiVRk+Yn3SQkM3UWzcXu07jZd6Pvem5Fob1fIxy9H3ejL1hklin4TL3+PXS6aT6vwGODBkjJnlyxjix4mOBTiMvRNMqvRfov0P0P5d+vGvg8b/AHkSv5dl6Iji3kY8iKFlTO3o/wDizu/ubuRNIWRG74oS2ttydi5dpkVxwizcKRHJ8eOaRjntnlcZYmxSPMFITN3Nl7RcmWEzfxkSnilI747LF2ui7LNxGRuL53mNOUopOM7meXGJso5rZxHDy8VKTVfejtpji3CU435rHcikdjuU0XwXzYyT0Y3ReljfCO52HotGyy9Xo/Tyjp88unyeEzwoz9KpY8snjy5Mvm5JT4eaMcH5jLjlB8248bRx2ikPj5F0ff8A18f5PG/3n5K9EWSScUfeyy9Lo37lLW9OwmIuOlllinRussrT7JikbtF+XHRhyCxF7RK0xSFM3cqYp2edQp0N8edtG+bHQ9bGxMiSZy2savYoxxyRObguZtY5SIQW+/i8rZFzockoPltxvLtQ8m0eRtVylxuFdrHuOESno5cW2bqL0tV3T50v0t8NlnZa/cen20sb0utOi8Qn0c34lk646jrcmRkX8WL4pZMzSnJzZBbyWO0ri5cvt6e/qf8ArY/p+N/vK5Wn20i6cpbmWX6LL9MR6XbsTEInk8ySY9GmjvpZfP3sWm4sRGW0bLN1EGr32SSbl3NxuExSNwpkGKVxcXJ6dm2XpXFcxjxGFk8W11QhqlAveoYNo5RKSjt2rLnZubN243bVbbll82KRRu5KsQ3FFn5S/hnInIfBRYx8uyyz7lifqaHxq/k/YjIW7IYMDlPruiXTp5IxfSxeeeSa3dP00sqyry5NtnLHFjgyrHEcR8fIr/Vx/T8b/eV85F6XotEyyzuXRZYmcFjZZJxl6LLE6L0izdRuLIz4LtebQpG/dOcXF3pZZuEyNtwdCyeZgUG5uI3WjZyI4Im9I8wi1uxU1LFuIwihqicso8nO+hZrJ5R5EoSzqbli5UBwVq9Ix3nlxibknfCtj+F8RfDJuKetm7ncNnfRPSy+LEXel6X6Pvper0vXHlcDwHKsT8QcOsxZOj2OEJYDN0c/J8H6Zzl1eDEuolhrA8UqjBkpqnGtJy1u9HrX+tj/ACeN/vP21r5S9KL1stxd6ovVaI7F6fZMs+yL17rzKN1xhmqFpRlJSU7L1ssiyzzKMeXZFZmZHbsaKLNxLg3FnYWWnilbmoYibeSWTF8GHqVhi8jzTmmTVEsu9RySJd0rFGicdpCJtoipbcnwPJ+VK3+UaSeVKOScqO8fyl2t43z2GNiRKK07jYxd6t/e+TuMvjR+h636Fyun6ieAwOOTB4gvM63HKOz3leVizYl0vVYo5Y5sfOKc4m+UZfnFB04csYzsjvp3LO/+mhmP6f8A/8QAKBEAAgECBQQDAQEBAQAAAAAAAAERAhASICEwMRNAYHAyUFFBA2Ei/9oACAEDAQE/AafivWdPxXrOn4r1nT8V6zp4XrOnhes6fivWdPxXrOn4r1nT8V6zp+K9Z08Lt49OU8L1nT8V6zp+K9Z08L1nT8V6zp+K9GRbS2hoQR9BT8V6JiyyLIvoKfivRLy8/S0/FeiX9VT8V6Jear6Sn4r0S8z+kp+K9EvjMx9ot+n4rzeGQQQRvPM+1W/Twu3jyqNh5n2q36fivOedj/mfCYSGQ8j7VbUEGhJLKfivOUPLDMLMLP8AhhMKIWaSbaMqSSKUmjCyGQ86Ss1JhMLMLMJhIRh/CIywzCyEaE5qfivD4ZDFRUzBV+HSqF/i/wCnRR0kdJHTR00P/P8ADpHSOkdI6R0zpnSOmdM6Z02dNmCowtdguTCzCYV2dXBRxkk0IRhRCNNySbTt08LwOGYWYKvwwVfh06jp1HRYv8V/TBT+GFfnf6GBHTOmzAzCzXIk2YGYCEPZ/u7VwUcfR0/FfcQzp1fh0qjos6P/AE6KOlSYKTCiF9jCMKMKWV9tVwUcfR08L6aCCGQyGQyGQyGQQyLKip/wX+LF/ijBT+EL88CfbVcFHH0dPxXYpNkMwsw1fhgZ02dNnTOn/wBOmjAjBSYKTDT+GGn8NDQ07+CPDXwUcfR0xCNDQ0tpfQ0NDQ0NCbzaft4tBHgT4KO+bFraSSnj62bT9HBBBH3TKd+bSYiSSTEYhu2IxGIxQTJJLvTwNwY0ck2nxSCCCCPsWUZsRiJJZJNpObTuySTkXBXbFA3JiYmYxVE+gpJJtMlOhN52JJJ2ZJ2JvQ9CrV5nenX0HN128EWwipOmYTCOmDDI4WhhKR7KcGPtZ8wWeLwzCzDJ0zAYB6Chj50P4Qv6f+SUSiUSOpSYzqFWpqjEKsbRItyl+ET9fOzBBBAjQgg0HaBIbFUSKoxGI5HqccCf6TBJJiMRJNnnjdQn4NE/bO8EGtqR2mB5Gx2dpyuMsHFpvPZ02mCTEST5zN5FdjFedqbMkkknuKSYG5ySJnPms5ovFos7Rac03nKrvuFdZpJ8knYknJOaB3k0ySSSSTbTIzQ0twTeLPfjZWZ+TySTbjMryc5nleRkC2XeLQRZEi43IzJEXS8oe/BFpzQQQPfRoNHGSewTulI1ZPIrt+czmiRoaIIItF52HdDyrNGfmyOSBZpyryV51lnLJJNpuxIga7ZMnaWTi0k+XzkRBGV2kbG7zaSSSScjRBG1NptNp30rcEkk+JySSTvQQRbns5J2P5abznd2RvrMsqJyp2Vp8fkm05Wu8m9I3lfZIgjYVn4K/p5tJJJyQYRUmAdJhurvtZJHmjdXjcfQtWTJJV4HvvbkTJyPem6JyT2q8hkSkasmTeru+CRbEbKeVdgvKpJkiCRVEj7xu8k9guyjJSpGtbLZXjqqtBMXwkDX0cbU3kW7yO9Lge3A/HaHqVcaGonI9DEMeWe6knem0k78EeWUuUNGEZxaCDgZNlruvI9uc8C7BCpkS3pvO4vFKXDFrZ8kySTZ2ggagkf0S3kPYkeT+7Mk+PU14RVJoqqsuSkbG5stR02d3svt0fy/8uh3nJO89cvPkaZyU0yOiCUinWyRwTZoi0bPPbRZdms8k3kZJo/JKXB/mNSYBacFVP8ASgqQ6SCCSLPPHextLa4yLIs6yLJP20k9o9yipq1a/wDQibNJjQjU5IIJy825J7f/xAArEQACAQIEBQQDAQEBAAAAAAAAARECEAMSIDATITEyQEFQUXAiYGFCBBT/2gAIAQIBAT8BxO9/WeJ3v6ykxO9/WeJ3v6zxO9/WeJ3v6zxO9/WeJ3v6zxO9/WeJ3v8AV3+uYne/rPE7340/TuJ3v6zxO9/Vk68Tvf1nid7+s8Tvf1nid7+jWo0x6+bGjE739ErQufLQkNz7Did7+iVp7rIfx7Fid7+iVp6GV19o/wAeXseJ3v6JWr/m9TF737Hid7+iVq/53zgxHNT8Sd/E739Errqwe8q6+J67+J3vy5/bl11YPeVdz8R7+J3vxZ2p1z+pTboLVNp1LVhd6K+5+I9/E73+8MSnpsf0/tlpSZOnD70V9z8R7XU4bFg/IsKkyoxO9/uUa8Pk9Uk2y/inbmQRJF4tCMqMph0/kjFTz7SUipga+CHeGZajKOmBp6srFhsWEjIkRpxO9/p0olGZfI66aTiU/JxqB469DjM4zONUcWo4zFjfJxv4cb+HF/hxf4cX+HF/hxTi/wAOMcU4pxUcWkz0mZHLfXUkk52jR/nS+mxh9xi914MqMplIZlMolG3lRlRkRlW3id7/AEKUZl8men5OJR8nFo+TjUfJx6B/9C9EP/pfojiV/Jnq+Tr50sz1I4pxEZ6TNSStDqSM5nZLMLuH12P86X0v/dOH3Ixe72PE737xmSONQvUf/RQf+mk/9P8AD/01HHrOLX8mer5JfuMszszN6cLuH12P8aX0V/TTR3Ixe72PE737NJKMyMyJRKMyMyMyJRmRJI8Sleo8en0Hjv0Q8Wt+pmqfr+hYT/Iq67H+NL6K/pfpajuRjd3seJ3vwo0QzmQzmczmczn7HJJJPu2H3FXXY/xaSbPtV10snejuRjdfCnwa8GamcCo4FRwajhVHBqOFUcGo4LOEcI4RwkcNHDRw0ZEQlaCPdZtJJJPteH3FXXYXZpfbddLIYijqY3XzlS2NRbKQPr7KlJHMgVJA0QZSLJWj2CSSSSfZMPuK+7VNl2af83XS762p6oxtp6EpGrcMVA6DIKj5MhkKaYtkQqEjKjKmJQRJlV31EpMjGoMtotBBHlpaovH6Xh9xid2wuzT/AIvT0dkPqQUdxjW5mVkMVDZwzhCw/kyIyoyohGVERaNmNEEEaH1KOlokSgyoakyDoMuqfDagZTzFy/QYvBBBBBBBGzR3GJ3Xgggysys/zZIymQdP4wcMVBlRwzKkOlMSMqRUpIvGtkWjRGmCNiL1LmU8ls1eMylNkDpKVBMk6J/SIIIIRlRlRlFSkOmWZUZUQiCCNK2FZ+I9CZJJmHUjiIzjrKapHXAm6uZLGLps1KTIPluTrSHTIlF3+ixaCNtEiHo62QyI0TZaZs9ib5kjOjOjio4pn/hTzHKFMcyeY2/Q/IhkMhmVmRwcM4UFPI6mWDIKlrZnTWtmdjLykRSvX3RKSPIm8aI1u7FogjVJJJJmM5mKiWSSc2JHQkbnoUodEmUdBkFQLkLkzr1Gl6EEEGUykEbM7tRUtlD0SJSUqEevusx50aVo63jZlksliMo3BnM4srOhU+RS1IyJFoSFZWgR1I1ydSNUeBBX0sqZMrOGZDK7q06KVqndf6ErzbpsyTqfMg6ikkyoyIyoggfNEKyFFmQRtQRfKZSNEEeHUZJYlBF4KqZGrwRZUi/SJ1rVN4ulsNC0zpjT0JFbMSTZWnVNovGl3Xlsi8WSkS/QI258GCCNCtGmB2gi8SZbQQKzYrwOVogykGUykHPTLJZLOolefBnYkfO7GTJSo0PQ9t+8Rqi0EaosltwQRaCNCItA0dCdKd2IWp7KJtN5GMjYel1RqqZmJtU+R/SbJbL9+i6ItGxF14UEbEknUjVmJJFq6bLOZJ10R4DUi6WbgTm1Ss7Masqdlke8xoWhaJtInad1D1TogjcjSmSUsTJJ1RqjT1FtSN6edulmJwZip6WZduNp+5xoSOZzIlEM/JGbkKXadC2Z2FremLQQQQQQQRZCZJIn40EaY1tknW0EaJ3X7nF3rTJJEzNBnJm62FoZJOxFo0SKobJ0JWggi8EEEEEEEEWTESLZjxW7QQQRo6a5J8B3ftUD0zeCEZTIZDL/AEhikcwfkfkfkTUZqiWxVMVRI60jiUyZrVVQZxOdEanrgS1Roi8EEXRIronyqiNLRAyCNEePHtUEEGUykEEao2IRCMqMqIOGjhfBkcQZGVU1DkpqYnIqvTz65Eh6F4c7LXgwPfeqPIeuPEjZjZgggyp9TIkZfg4dTOdPUzMVbOKjioVaMxNn40EEGUU+HN50SSPwI1Mm07D2X5MXjaqGzMSTdWaYtEEeFBAn6EyNDoKsFlVDpJyqSmvMikV140EEaFvRdkW6aOvhvVBF41vS7O60rcjwssnDRw0ZSCLx5eUqqdPoKqbOkdLR+VIm2YflwQR4E6n4DtG++VmTCJkkfJCc70XemN6NmCPZHSh0xzRnlwIyCogp5eJO3BHgPwsw74mJlcCfKz2anCkprkqcdBueYhpsgak6DKWSJzd6+mqLwQR5LWvp5cFWFTU5JjkZ0nA1IrZxVCfuEDW4zo5FfFoziHoelqTEbiCinkOkyQRBFoHSNEDREXd1pagT5E3jTFo0MXiRtLyMSnlmMFqeZyHTBT+SHQIWpeTHmvRI7K3XYZl1O7RHpZqyIII1PoKbIgWw7IdlZaVpm0kk+VG21Jirhv8AEodXqU47bgpZyfS2YkmREW6HX2KfBZmgb0Rp9dMXiz0t6WrraUEbUDWh3nQ2TrgjYi6343aqVUoZiprkUtop5oVLS5EGVzIymqbSSTJAtjr7QxdY2IgWxD0QQRtMa2ovl2mRabNEWkdp0ogjTOrrpXlYmEq0PCycinDVmirkKkpUWfIVR1F7UxKN17CUD3IvFoIGRoggi8D3U9DOg3oSvFojbgjVG713mjkiuqEYeJmZlbK/xEiutLkU8xJKyZKJJJOvuT24uuW7F4IIFpggYyIeyyCLMkm0IgggggiCSSb9Cda1RtRtxsVUyf8ASuiRhzSxYk9BvN1KcRTlMepdEYdbyirmrmZkSiCfSyXvHXQyNcbcWashanaBqeY0LUtDQ0dbxJEIQiCLTZaVpi8EaXojYWhbldCq6jmeRhcqBrmZecjTzSUVNchMcdSE0dB1GbV08r//xABGEAABAgMEBgcFBAgEBwAAAAABAAIRITEDEBJxICIwMkFRBEBQYXOBsRMzcHKRQmCSoRQjNFJigsHRJENj4USDk6KywvD/2gAIAQEABj8Cfn8M35/DN+fwzfn8M35/DN+fwzfn8M35/DN+fwzfn8M35/DN+fwxlNcE/P4XyU53vz+FvLRqn5/CqSnfLRfn8J+a5bN+fwl5X0VdjVPz+BkC8F3ITKxWFi5wjCL9Vb1kzuwkofrbOsPd/wC698z/AKf+6/y7UfhT7J1laNczeIGID6LVtGk8o7fldTZV0X5/AlwHC6DhERElBrQ0dwR6VZiNmffMH/kg5pi0zBQj+8PW5tlY63SLSTRy71gGsaucauPNNxMa7WFRtOKoq7Guxfn8CbXO6Arfg/4W0Or/AKbuWVxtH+Q5nknW9v8AtFpX+Efu3DCeIM9OqqdlXbPz+BNqe/RdZvGJrpEL2HTrTDD3doftj+6HTHe4HuG/+3Yb8/gTa56XQv5v6LoXh9hvz+BNrirHhpdGtvsMJB810WzfvBnDqgaanbvz+BNppHxGrox/02+nVLLbuz++8RaRFFx/CVF2ID5Ct1/4Ct20/AsGF7TCMxtTpP8AnauiH/Sb6dUss9u/P77kQktbd53RKxvGty5aM1qxct0oAyJ5qWiIU5aVr8zfVdC8IdUs89u/P78RhEcQm2lridZuOEYaprjxEchpBYx/MFj4LE7eP5I6GHC/OCbBr6hStG/Ve8b9VW+2zb6rofybPWcBmtUh2WwZsZr9bbsb5p+Bj3EGXev1Ng1nzTUH22EcmSQ/Wv8AxJ+f35s8I1fajyVnik7CI6JLrVsuAKxe2GXFb5dkF0lrsX6M0A2bIUKlZvJRwWAHKJWphs8gji6Q/CUYWrwDycqz0IteQc01wt3xbSJQHtMbeTgraydZtAMJhdGshY4nMECSU0m1wk8CKL9os/xJjTaNxP3RGunbWTMIax0BJB1sYwEJJ7LXFiLoiAR9tZmznLDNe/8AyKH6+MeQWrjeeQCOGyfihxXurL80/wDSwGcsATXe1a0fxFNew4mmh0IutmNzcvfY/lCPsLAuPN5Rw4LIdwR9pbvcO92i3JPz+51VVbwQiarfC3lIErcW4t0LWAKkwLXbE9y3Ctwr3Z+q92fqvdn6r3f5r3Z+q92fqvd/mvdn6rccphwXEeS94FK0afNV27j/ABt9UyNpiJFGzXunRzWrYtGZRBtTDkJKBtHEZ6FpzwjRtAZhplfTRtMk28EEgihWrb2g/mXvcXzBHELN3kji6OMXcVIWY8kHYw0gQkE5zjFzpk7PCLV4A4RXvX/VftLxlJa9s9+btk3JOz+4dQt4LeC3gt5bykCVJq3it8qZ67VStHfVb+LNa1n9CpxaveBe9b9VJwOhF1oPJGAc7yWpZAZr3mH5US57nTFSmZbB3yaNrneLPRtMkOwhknZ9sTIW8FVUK3VQLgt5bxVT2jK0d9Vv4s17yA7tE5hWfyjYO+TRtvK9vy6NpkvPsJuSdn2NCIit4Kb2jzUnA5FVCqFvBbwW8FVQxBVum8KUXKTYZre+im4/cJ3krL5RsP8Al6Nt5XsyN0eHFRutMkc+wm5J2fUf11syy+YoMb0pmIosPSbIOFRiU+l2X4k1vt8UeLRILDF5b++GoytPwoxsbSKMeinug5S6L/3qXR2jzROGzhygv8sfypx9tXuosPt3KfSLT6rVt7QfzL9otPxKJtrQn5l7x8/4lDEfqo4iTmq7KqqdlVVvoqX1VVXtNysvl2A+TRtvK+zyNzgm5XWkf3U75uwhkukWT+jNfgtHNiHQ4r9ld+Ja3RTg7nTRxdGeGdxXubaPKSH+GtMPGaP+GtYeS1eiv83KfRBi+dGPRmGcpohllZ2Z/eE02Hs2w5NqvetZ8rV78fgCJ/SrSJX7XaeRU+lW341ie4vPNx2tbq300JGKmq9fqq307NerLLYM+TRtshfZRHA3FNyTFafKn59ZrowUlG5s+C6Z4z/XsbFxKiFEIRmoGqqoCqnRRUlVV6/VVupdVV7DtFZ5bCz+TRtflF9j53FMyTFa/KVa7WRUChdRZIl12pMqZXFSJgo1UqLkqonEplSJC3jc3JdM8Z/rfHTp1t0VDhoRadCHZVVW+imL6qvWLRWewsflOjafJfYedxTZ8E2dCrQ/wq0CqpOVFvBS1iqKbVqN+q/opGCh7Rb5Rg5TN1dOuzbkumeM/wBVC6SjpR6vEyR4JzeSaeCj29VVW8qqt3Nbq3VS6q3lVbwVVXStck2+q3lVRQkrE9ymVGKM5hRBTrRxhqrVmjzTCeCIAuwxELsJMoIwMFU7Gl1OrNyXTvGf69gGHBEGZURJBAfZ0o/cjldIn6reIW8VvqqLXGRQAMFvXVW9dAqRmg4nzU3EqujTYV6tIFUvkqIxkt4Xbqgm5Lpvjv8AXZGaCj1Ikp2CnO6ey5fcSIF/EnSjG6BvhMlU0J7Sm0lobwC961ACaAIWqJKAbNawipNP1VFRUUgowVLpXTXK5uS6d47/AF2kDs5aWFzcLUNeCwYo5dqSW+36ojqhQioQvqq34bqKl9dny2E1I3ViuMUcQkiBK+P5KQXJc1rCKopBTXcqKklyWGUFqlT0KbRuS6d47/XajnsDNQ0owUUJx2/LsaXFV6rW6uhLqM9Gqk+KrdAKYiowVFqiBUCq6yIUVPQrBVUutNyXTvHf67WNbweakFNVhdndBCKpO4rWEHd33DndLSmpbOKF0LoQVJ7KZUYqV8CSqOUYoAO/JVUyVJCVUdKfXG5Lp3jv9dsYeSnpNUeamYzUULsNUNhHsaHYXfsJ7OmwHPTige9HRPXW5Lp3jv8AXqwio3Gam6v3MrdXsg3R29NGq7lLZNyXTvHf69WnoUhD7o5dRl1OimqdgtyXTvHf69VhdD6qU8lEGaPZ/fce3u/Srpx6nLYtyXTvHf67Sa7lLQlowXJQBjsJXC6vYsEepxWSotaKkSoXhcroiid9ewpdjNyXTvHf67Ot07ip9Zr2BHqtVWBWHgioY6qKoqGMFulUiEYyQAfVFocCoRgboqH3EbkuneO/12sdhLbVunsY9bI6lQKBYFSC3it5c1uqkkYBUIumJqQUk2UFK/uRuku/YRhtYx67DbtyXTvHf69m17MF1VW+l0nKTr4YQVH2YX7OFAsX2lrTapRQrFQDyAjG1UBajzRjrR5LE78kXAat36thcsTmQCiVSioiiO2G5Lp3jv8AXsTlfDZxun2NP8lK7nfTYT2FVUreKjFQbaFqHtGC0zWJzIDkEYtksJJEeCAxCiJEA4oipWOEW9fEVLqzcl07x3+v3ZkioaFY6NeqVWofojrFAuWrEvNQaKLYMHJYYrVKxKTUYtPXc13dSbkuneM/17GpsQgo3xu5bSfVyYCKLiYRQW4e8hExUlALndG0GPuWqMI5dX5qB1Qg+InyKEoIoxaIJrHtxd44J2qGO4I2b98Vgh6KnZzcl03x3+vZcADFQa0k9ymoXZXBRFFCqIWHhdOm1j1WUVD1VFrGXJUvmv7aPK6vU5LWQBtQzvKMJzW75ppITXNtPZuI1ophjrA15p+qMXenGk6dmtyXTvHf69eHHYeUUWhwcOYWGEHd6GJ2pHWMNZEWFIw9rBPLWuNo2TXNNFb+0xWdq1sgJIOE/wC6mDO+ChBZqKio89vC43x29VKqMVMKmhXTr1eqwukI8F7RuuxxP0uaGlwPGa1TRtXdnNyXTvHf69UaeehaOiJBQGiL+V+EEA96Y84bOUINMZ808W2pFkGOensfYttXcDH0UX4scyY8UHQ1uSgXHDyQLxGW6TwTX4cLOIJqsFriOtug0UZlo+0THyWJrzihDD3qMYtvP5IlRvgqyWqVPQOy5dWjwvio38+tCaLA7Ew8F7QNr/8AFF4Egpt1TKPZzcl07x3+vUxGiDXUGg+US5V0ctGMPqg8hsOA5J1DGQQDxiDfRNdQtMu5ElushldXILDii0yxqDZu4IWL5zjHknCoE8TUPaYcLufBODTKNdCV9bo0KDfVSWq+fK49+0/qoKVOowUNHkpV67Z2BbjaTD6posQWBgG6hxG9NNBkF3Gihw0JdjtyXTvHf69gzuiXgQ/NYd71RleOd0VFADzUQVjdx4BS4qdmHDvWq3WjwRxNhCWxDofVRILO+KbhdLmiOOke7TgUCpc01d2hC6MYrWUBS4xVLjxUwjo8ro6FeshzDhcOIULZxfybFAWLPs4ELQ2hDgJhAzMVrgjO6lxn2O3JdO8d/r1ExMOM1M6BlIim05ruURJDjoEaWJCM8ysQwxaKGcUw/b49+jHjotdCIU6ckXAQI9Lq7SkkYTw1CwtFUGxidEmMlK6oXPvUVTvXFp5QVYbCPBSpd37GmnTaB7aqytNUvJm2MYIlzniU2rEZhsgiXEkoCK9lvRg4lSBUxC6Y7FbkuneO/wBdvEV5bCmxhDYC7vuheZqiwymq4Qed3Id+mV3qJkjDiNqIlTKhCHetWBJ4qUVMr7KgsQFVUrncYmajGKEVCJ0IL+yMo6Nb6zUzw63EQd3FG1x4CeC1uAww7ru5TUICV3JQ4Kiou/sJuS6d47/VHSio9Vj6aE9hPTkpiSGHgnHECp7Cd0h9diNCMbooD2eHvUVRREyomId3Ki/ugIKEFXyUwGz+yhUqaN0AgF6KIXeo8kJ6fffTrQlHimymQpICohFQHBFwBhzR4jQj2C3JdO8d/r2DNSENrCC5XA1cLomJipjYnmJR2nEqGEzXFfud6B3lI6q3oeV8EIiAKABl3VRnf/W6UUJqApfCMlVUKlfGGl3Xnq9Va2rmRkoywl2thRxGDj+aJY2fejakOaTQQqsdq7DZUgnCJDY8lAVioicFRQUeFw683JdO8d/r2jFQIiOSooTjmh9di9sJFQXnspJsSYHkoAHEouKxFxgtzEc0Y8VzPeooIASULo6EYyKwrFcYxuLRMAwndFeUdhK6N56tAHVNQiHtj9pUwx5IjBQxjGcFgg7W/iTrN1mTxBBXt6Ay+iBBMMMUWiE6qEZKajGKMJdfbkv/xAArEAADAAICAgEDAwQDAQAAAAAAAREhMRBBUWFxIIGRMKGxQMHR8FDh8WD/2gAIAQEAAT8h/df5EIQhcrhIXCROELlcIXC/QX/Nv6GP9R8Plj/Wv0v+sf8AQaD91/kSEQQkJCEiCELhcJC5XHfCF/8AEv6HwyjfFGxsvN5Yy/U/6Z/1b4fGg/cRcLkhCELhcoXK5XC/+Hv0tl5f0MY+WP8AVnEIQhOIT9af1L4bGUH7j/IuELAnwhcLhCFwhcLhC4X/AMG/ofD+h/Q/oY0QhBohCcQn9Pfrv9O+XxoP3X+RC4TFwhCExPhMT4TLymXilKJ//Bvh/U/of0v6WX9WlyX9O/oz+r0H7v8AyITELgiiYnwmJiELhC+hcLhfoL/nWP6W+WxvmlGylLwvNL+lSl4v0Upf159E/opxoP3/APkSEhISEhIgkJCEuEIXK5XK4X/wr4fL+t/Ux/1M/W3/AEb+rRH7r/IhCEIQuEIXCYmJ8JiLwnwuUJ/84/pfDH9L5fL4f0Pl8v8A4Tv+mYzQfuv8iEIohcoQhcIQuVyuVwv+cf0vfDH9L5f0v6H9D/qX/R6+ifVCE+rQfvv8iFyhcrhMXKFwvoXK5X/wTHy3w+X9L+h/W/6GcwhCDRCEIQnEIQhCE+hohP1JxDQfvv8AIilKITKUTExMomUTKJ8Uohcr6L/8Cxj4f0v6X9L4a5g0QhOIQhCEIQn0T9ef075ZoP33+RCE+ELhPlMomJ8JlKUonwTEylExPhf8w/0JzOZ9DJyx/qMf9Y/03xPohPpnLK6BJD9//kT4TExCZS8LiiZRMpSlE+FyhfSv+Xf6DY/pf0v6GvohCEIQhCEIQaIT6sGP17/UoSzgbaPuzLYTBoP3P+RMXCF9FExFKJiE+VyhC4XK/wDhH9D/AEGN/TRv67+k/wBWE4hOJzCEIQhCEIQnCEIQaL2/R9gJFnb8vhC2xvQvuyN/afuf8iYmXhCF9aFwil5QmJ8LlfShf84+H9D5f0sn0wnCEIQaIQhBkJxCEIQhCEIQhCE5nMJzOJ9c+hjaWzPSlvb7ISaKDaW3DPSlNuekJdFxoP33+eELlMQhcLhC4QhcLlcQS5S5XC/5l/qvh/Q/0Wvpn/Evhr1l6MthKs7+RtLuGelSNtz4JX06BPy/5EEVwILhXGuBBIJBJEQhC4X0IXC+pf8ANvlj+t8P6X/ymhr1n4PiHtn5H/0Ct6/It7/ASIhOGPGyeqz4EYGR+6/yIQuEIQvqQvrT+hP6F/zr+l/ov6n+k/6Jn+4IyIyFMzkia2n3+xtv1H7mobG5NnZ/9sH/ANsf+4hbKebWlaGk+MD/AB9UJ9TaW8HqmzLtB+Tp6MZ9pEd1/Iklr6Gxr8/BT0p8lPf4Erq/POiP3H+RCELhC+lCfFFwmIonwnwnwnyhcL/kn+g/pf0MfFH9N/XnMIQhCEIQhRivHUQe0Nw+T0Z6Q/t9nvD2u/KE2FYNNG5T/CKvIlWWWtJ2/pCw9tfZHbGiZ93f6LRdklvUMvy/YrwRXf4Ed5+TDS4nDR2eibMuki+/wPUQhBog0aI/ff5FyhC+lcLhC4XK+pCFwvpX1r/lX9L+l/TP0IQn9BetTXhrSnS2/ZnwNp7QtLvv3pn8nQp5rM6yWE76k9saTPr66k+P5PkxJIqs9GfYNuz5I+SKH2o834ojtn3PUQulw08k+Sf9R8GXwJ5JF+RHefkk5fEH9K0hfzf5EuELhLlIXKEJfUuF9K/+DfDX0P8ATf6U+mEJxCcziUDqe5vRIQ3oUDSo7E2C0Tfyzp2KRvKd+X+eho4PQeojwQiGvgnwSSSR4J8IjwTmfoQnDJytIT83+eELhcrhcJi5X6C4XC/RX/GX+if9JSlL9V/QbhD/AGf24bh+zhi1ixjwQl/SXi/S/pZohPyf5EhEIIQhL6F9a4QuF9C/RX/J0peaUpSlKNl4pS80YpS8UpeSlKXg2UpSlKXmj8D+SFju6aPQSLw2JSlW7mxP4JmxWrvK/pHGfoE+hogmFk/cf5ELhCXCQuUhInCF+ihcIX03/i7+jS/RSlKXil5v6j5v0Uv6lhl+kSFhbsom3y3DL9EhZnj+4e5P4n9Jmostp/pwhBLCP3MnOPrpSl4UvFKUpeKUpSlKUTKUvNL+jS/1F/Sv00peaNl4pS8X6H+o8CXoMcNJvJbt/wDbwbzRK/8ASU1/oehAm8zmwt3LJjT+/wB/ohCDwZfDRG/RgjJ+I29GiN+hcIW9X8x7K/gfRCDRCEIQhOIQhCCEhCEJyQnCEIJYR+4/yUTEyiZSlKUpeSl4LgvJS8lKUpS8KUomUpSlL/zr5g19M+icPGduwbg10T9emKlse9HU7JEDLApWhLndEi3EHHEUcn+B0zqQJW5LhONrQlLCtNLBgQhCFPU4W3+sITmEIQhOEJwhCEIYCWVUQhCEIQnCcikWR/zf5KJlE+KUonxeL9CZfovN5XCFwil/49/pz+ghPphOJxa8xjzCBE1uSP8AwdlagZXwT0NuhVljzNw6z9Ha8mUqyxOypqXg8PA1P2dI+GBppS35Bahfo/yXDa1qaO9xYiciRv0+IU7f8Qf8P+7JwhCEIQhD9wFBbUi7akIQhCcML3fQtLMfUCEIsyS8sRp09LJmKHyNJL3FU9m1kFj4+OtsbS7C/m/yQRCfQiCQv019C+tcIX6S5v61L/VP9KEINE+mEJwhOYQhDaRHfgyCtA8Y4Y64hK2ezX+W6H+BJoT6J/sLUaXlyLauQexn3dyIyRO1xtr7n/I3qIjScn4FE4NMyQVbNnXk0XdstfJ7IIoMvk7k/JFUR5xa97LiNDyjiBW2YoGrmQ0JvGldRQ17R8CEJwhByjh2RbFoIhlfXMdIWmIJsE9jWu3+3gZEQsY2Mt+kf5ELfVhKbi/2fJqiTOfzRoC5jA58CkKdRp8QZLW0l7HZO9B3RvD2IU6ZAhUjuXvf5Zn1tpk/AzfsYwx/wBfzf5EIJEIThCEITiE4TiE+kv0Fwv1F/WXhudnoHrfk/wDQHcOUwNX+ca7k/sIDGFhE/kfifkjwkxpfCwNrB+WPQm+Rj/2h/wDZfRhGPf5AY/LHmAv+2Gf4Qa2/mCXV88XBP0j+/EITmE4ThCEHTbp4d6EM9IQWeaohBHXljFczVPpHq/1weVkzcEbFWZLtCfuManwQ4Y5XBeptHYTcLpj9xUjTJHydv/VG+3f5O/Jmmi6Y9Db8IxMY7cLGD1dWILW/RxRdj/f/AHKfARYsl++o7YsCG3C+hrkucJDb8DZBs1syuxOwSSPEPObn8xZTVSkf+wSbryMZvbZHyTZIQg0J+AL+WQn0CEIQnEITmCRPohCCROIQhOITiEIT6p/SNF2hp/zDX/kGj/Mf+sNXUR/6C7EYTwvy2NHivgb/APKbEfy+YNfU2NjKXh8Ph8FKN8KjHCzEyIMP3Hjz1pBFt+Q/lsqdLfKZqgftgPli3lFUsmxRRdTYrcjy9HZ36JBqpdsg9vr/AAMHVH4DsOhpLZIzR9P5KcGPBsS/C/g29DRt4wz2orfRihpiEpb11+5n8jGXga7G4N68FbZaUTc+gkzTgzL4lHkMYzJ5PXFntcTGiYJxm0aP2I/NvoEIQhCcIQhCEJ9M/RX139G/TeaaMfLP7JCXZ/CH0sGnX5s6ShjtPsNdvsNn+Ybd/mKfZeL+jSlGxvmjY39DGPhjHyxjHzfY+L9AU9wSY4a4+xo5dZ3WJUcL5FH+wNDGg/gGGo+3FJ5P8xh+XHKJj9/wNcDFILNf2MSEiVYZpoT0nT6cS9Eo8vRgINiQ1wynRoa0dcRH7DWBLw1kYkWB4FgiMGaGhjydB0P3D60iE+icT+l0SltQRmU2k3scpofhspfcBUx4f+0f+0f+of8AoGdLK+qLxvyMiMa2qJmkI8n8UHTSfgFWP5DwX4D2V9yeWJFWzSFnP0Mf615Y/oox8sfLGNDHwxrhoY/obHBaUr5afIz+c/kW/wBLBXrk9h4j6jfB6d/3GCGuNP0YH/WOLKRH+2D0CkcghEuujQS4Tn6XH+4ydweMEJBqrhMEiOw84I/uaXfklOtiehVrZ/Ik7ki7wMspkZa8GQ9hrHCXkYeCC9nQ/cCcwhBL6J9SQ1D1hGUzIk6qPbwIuBHfsEZFryx/IJmNXQvgfacxTZedlmkjwlHUULs/B94HZ/f/AOg2PyzscJfqmP3HeTR4QQqerSfAWGl5SSf5hDTk+JdynsJ+X+WewoWZFd2rCkmn4oqTeQYpq2b9sTvseac4L2ExCF7CeRq7L7i/7gTE3kTeRN5Ym/JX5K/PGgbPa/Ikdj2HwHoC8ivCxewuPUPSI88v6H9T+h8sY+GuGNEGicNDQww0NEO+KPHNEzfDKYe1/JX4g+A/UYQsJD7t/eNH7I9w8/I4J68fxHEiNLwE/A8oUZgvgMJ5X3HtuGTMD/1DUcYuR0/ZjsyoYxGiLrYi7RuYGaFloydmBE/ZFF7DTt7HYUVsR+B2TYvgyzMg8PXBmG+H4EKPiy5EyF3fj/4L0c47AyqMw0t0Wbo9P8jU5OTS/YeEZOHaZavfUD9pfD+DZ3Z5VF0ht3aoy/JlR7MDFRFdJyaX+h8HYOWrj8G3/CCDKXyPmroZazsDycNp8DNNNCvgVtQs6F8rgMm98ArbYp9Mohto+KF2sGLSYwVRoNNNokKCgkKChhdjIk1UKJGkZrMk9sasSmRgq5EIICpSjY2N80vNNGyEgfELtS4k3aaH5DSvh8v6GThjQ1waIQg0NDQx8Mg0xpkGuL6GXGvoVFwn7P8AJnwb4LLH5RroMUfLhfBMF4S7IU1/YSGKd9H4hjujUFKOJ2rySzYoR5aNKZG6EL7Ub+KNRZG35H94iDVcfCR4Mq9G3oj+3EwbfJUyTI0tDU6JXFscW8GhPwJCY2I2Yba7GtZaPRkP8ZC1hJeWag07Ml/6WQRYj8DQ0FAlSPJI+EI7gakPjIg4g3nQkXgSsq2JaR1Sf9ZXXDoyxBfcJJb4WXjhIFC4wyCjwQSWNPYhU0MkMNNk2gP+I/UGxJeSHSqW2bzhFwTkPKExi/sZeeDzhRStFJVE5Kny84UXF4f0MvFKS7Egr+SewneuF6Indr6WPhkIQhBonDMjGNUaGQnE4ZcIThf2v5Hp/wBZEhpEeCX0PkJe9jNDxGsi6fyMFffA4H7f+Bn7Cfsstj6CH8r/AIE9D+0YpPtMYnqMcDyDXXDD3wZZ0eRIltmxsiXiDQtpdD1i/gpb/hlKXL68ERu2GqnpEWkLuFjS8mJVPuTDewa1EL7Xyg1r9YyQzYpI9GOt/BGkVUyfZn7H7IA9v8g2Gf2hj/uZipUb0Jg0NbjwXFFgS4LE+cIbPpxIqLPYKmRJvhPyIJAl5MUSKwy9CcPCio+BDRofyKEHpsR+MFrIll72ZO6gsMRBI0IE7MjDZSGbcHkIZsUQTg14UTxwnwalChUj24pMNm1DzlLxeaUf0soxjG+F3glBL7TPQhef7xdwj5T2FepfSltNFT4hBhBohBoa4aeyEIQhIQnGXwr+Snov8l5nBhox4oD8zLklj2yNPchItDT2bCx/0MmLxtVryYkjnkLhJ83oQkSyxl3cPhCxtEhlabVEN2LyZNXgTK5IlB6W74GJq7Ni2p4Fvbe0OraMZX9wQkU/WxGqP5E2tTjExSxP5Kn0N+w86E2vknoPoMOx5iibH9xUIXCZHgYaUb8Qyy/+0Qs7DY1HThJ7TGbhuIhD2jGeyUQ92I/mbmQoWBWQudEFQimGKiGhLMFPGD70SJeOJU0KqJUsFYx5E889qvYpJPdMU6r0Y9uQjfORoyVJi6jFAwQrE2a65bFwTGF9CGGEbGboyYtuCesCYny/onE5hOGhrhvSHjh4RodPuNl4Y2WtMhr7fkl2IP7yXR/Yr2vwQ5SCcJbnD5Ogc/aLMU6DdqfkyRU+RaiF8JfyfIy74hPYz/R2MsrjrEPsbS7wYCm0knk3ifkoLq9CIrIhXq0J1DGv8lylewVLfKMaVwL/ALjHVJZ6a6G9x8xiAfRtTQzLTvBQmml7Q31T5Iy2rwOusb9jbrjG3oY7CV4ZKwyGoYKCS4p4WY9J/I08Dwoa0x8klaU80bNn7h7rohINkwx6FMopG8ofyTowh32PDZfTGd2hdb6/mj2MXM4aEQhgOzawoSZiCa8q4kE4oMWRBKhHs8gh5CsGQcK20YtuiFfYLu4rlowDKiNV/gzevJmRmC+TwDfRCHkgoYguGI3Fci4T5QxvmicaNiZc1+j0Mo2zsqG+GVCHx4Byex6RghjbKDsiG6zZCo0HHVSENiYKdDWghjm3ZR4GlvX3GlG4Jh4qH3a9C8jvyRygwq4+4MElssxBc2xTCXXZGIVFG3yLFmvVY7Nz7RDTbqHkbbqFK7A6bhRjBCuj91AzLYTM37JYSwKwjpcpsdSHlBi6ECnYoQl+rTE30OI6IHXgS6Eh8h90J2X7mnLCpPJCDiElTFHYm/hFx2Zehq2aWuG2mUJTexsvIXQKp5bfiFkj+6F2QldB5ZF0fJi/nZvmXdGexvD0If7mYhkzw+N89iGWX2CyrL7ExaI4ZD2/YipDMuhSS0KnwaUX3kWewufXGyokMa1IVa3H7H5F4UhSGZE/wN9yinXgtp/YTYVr9iVJCCXYlkSsSOgh7i/WH7jEuzzFB0hRspRsvGTI0z7nWyXvk/ceQ54PAs8Eg2xPIw4LwR9kV74o5oSZE9j2hq/gautGyfrgEpH2NqeCOTJjHMn+4EMk0QLaLBHlSpddDUQV6MTa0MvAhnaIRZG+ACy28HDMLwNpjJdvQmxb4FfRkdkNsT4Y65cYyuvAk7H5MSNaGl7PZYiTIqVofIZ6CbQrDN9G9bH6i0qLAViihWgTei+Tob7EVwdv5jFmfYFTGe2h4JGBc/YoQ/IwTPkKydArcp7Y1uv45Fp1+CI0fgmVtj85FoJ35PBk/Z2TEhP5NR1PTE1dujtnof6zzL9KNBb40jAzv7DFX/QkRfY42ZK6F4IUUY6W+JomEO6Cn0Xzs1gzBE90YpJR6XktrjfwJkSvQrEsCL7mTEIYDxIWnHzIsimEpv8ARUXIiCXLc+hslTNmTLHQwyEGyoZS0nFQofHNN+TB0+RpAT7aHTG80UaZGhOkU1ngGvYhkLfYY+jyjeR2leE968GwZQrBY9PmDbXX8DQx46EJRyl4omrdopGmPV11sXYyonRHGCNLcRjy9DRLLMaleS6tQcpYy3JNN+yg/Bu+BIhm+D7cjD2KzxkzLBRpL8i42x3NY3h0jMuyEWRmbur7Eyxk/KJnVD0JJjKwPkKM8LyW7V3oaejqDjpJPbpg6NjPRLoWp4QcEht9s2J0U3nZCgl+Y/JQGye/ogUqDifMJU/4Ny8BhS6Eq4yVkf5InQMxhdGfgmBpEND8MP8AaefLKJi4ZBCQ2K3roRNVdCa1GyNvRtWtCa4SFQ1iqUo2BQ0PMnmGNvKpS9D82x+bMvgYp0aum4xwZRmGy+RIoxPtwlnB4dkSbMlCGkkecsPuBgSY39nFuLBCCFyLhGhDf01iTEwtfoDxGFQ8uLDbyMuuMmYmntBwfRqF55GEMbSH4Da4cmIZfJVc4EjIg9Y3UHl8GPBZGqI6CUwDR3sQ8tnY5bTJeDds1Z3tESlu/Ayjr7HdhDseup0Wx6xYGm56JO2hwngrOx4UT77Hk2XsM6RQdaDYyPprsgm1ckC9hXkHwXtvH4E6yjaTwU2iaqV1RK5u/CENp+0lJxPa0Nfb2eTrCo+RNwzU0fsbT+1LLajG8j9iVPZ5GGc0MsVFaPRKM8SxEWWNj9RU0hsDFPAjZmtnS+DKYFAwg2oQJqkd4L5uh/tPPhGiC4I2IyGjCOUiTe2TZUZNPR6S3ZsF7EIkyd4OqUXlDLVNhHHanQ+KeBC7WZlG+BpbiLjJVK5GySu3wzI32L9z4iRTRTYqwJXAlxudfgwqT1oToT2fmJCDLoSE9CFyQQhc0f0LZehPhRMQ2WC9jGiMbcVI0bmx7KNoxTsbNxlBGI/cV1E0Y61hm07sdDyvY3Q2v9xMDr+wGrb7Ri6xrb8+RO1oec7Kda/A08GJfsJ8A5hQbb6H1WeRdK+5mAnOT4IXAeGst+jLJUVrzD8J/wBge9LDExVKjfDaHjsdu2yjYH7E7CCboU7Y173cUc9t1UOqlzgbCR5EHD32iFFPgfbvpFtvoysvyN1LaNsa1GwNjMVGfkIEo6DKaHfoqaR2JGxoaZMDbgmc6Li9E+BoxGzISjRjeDodU6Q2amI62aGKMtPQ/wBp58LHCKdCyIXEEQXMXkUg1xl5LRsmqpa8FNaUN322uzIkkNnBPouiGdEdNrsRo+w3G42xuI5kyHNp1ro/YnwaLw0eht6N6Fc9BDzWR3nqmi8M1L/AqZF/JDYyvngTT2IohPkT4peGXilLkTLwuKKCjjFct6HwwhsoKMYo3y7g4mIeWuFZ8XtUMuJkauKDIMTXyGPOmJzA1wexRfAbJ/I+37Cx2YiuSQX/ANDQoFvwUbSyZCmhHUl0OJTXYrtYF59CdLUUZ9jep0OaE0RDbkrK9xvW0PtoxmDvfk1bhKhFMf3FUM+wxPoaaKbGnWCMj7h4EH60dPZPkPI4YcvAmwaHS19xWOZkHH2FuW/A9lGh5+h46Ho7KNIboayl4VKMaqJlkOGykEqIvsD/AGnn9CGLYvwaZ6INI0yTN/RfA3UegnXxk4X46NqZTTH4W8sp6zcibdNDqVeiuSuEIDCdZgUxYw0ef2NvRFwImsrJ/AwsQ0F1GwPOhvRmhGBcLhnwTKUTLyUo2bcGp54Q2N5ka0PKxEngVFBucORRi36KoYwwYzyH3Cria0XSUMfnwZcCGl9xdOps0kKo/wAjRNbHU7+DYaHWkarN3RYp6Q2/gUL5G19eB5f2QysCswXgrPQ1Y0OtumSMdaHjeiK10PsZF0o2muxmjXCy4QvtHMkTdTGf5kNi1gm+SEkwNn5H2AyUK0JCRgGiWM8OZgSMDJUlsDcbIYy2JkfQ19wmk8IZDBiyiBW7eBdh/YPoD3M84MmeEHpwnBH9gf7jzJyjBROF8C9HgknfGxseCCwhKzF7Fc3vBK3RWzCZs3DRmrdKfI/2xRkXDAgti1gRehOuF8kf7javR4QwJTJ8Bgs8GsdFHdWBvsX9jTgwngTExCEJl4Uo2XJS830ZhDZLwU4a6Efgck155GJ8ioZWcEDKxeC3YkexMDGPRkFUxOo2bHYtmGi/MiN/ydPnQvrA6hJMYYip2+SL19hTXQePEZU/Y3/oz+5gMNCCFmiX2QN4xkQ8DBjtHXs8LHgNlaFi2XhqmYCxtzV9joxHHZJHwW6v8DEVRV9jIwTNSGWPBD6yKzHGH+CJo8g5VErJBpeRVpopM2JTocImNEnoiZyQ7gcejRM9j70yU9RqxKjQXtCu0SnYmL1dDL/UzFCpG3KECwbgmL0zyneF7JkTon4Gt2NUvPaJTzwRUz7CwkFJPA/bAxrD23cCjoX5GAng9hY9mTFvwRhMXZD5F7Qz2RuDoVLyJgJDNoT8jYGQwuhd8mExvleW8mnDQ6E/YgwlXoRgyRKMaG+RieRCIhIuVbVHqHAp2NngwseaNBqQ0Me4v5GyGjA4agoQnQeFw9jmd/A509McmogsDNKzGjB2NnYm8FGPwPNEUzHexqM0N6z9uLTsLJc+zMmexfDKoyfkZgYVDc+Roqyja9DxIY1BgxI0StuIW4t9sxmesFlclJf3KHAr22xLehtfQT0Ssi4EP/Bcm3DSg0dPYp8htjKei3ZcieIN0SskVeDSM+x4RohqVbH5JNsbSD0WZOq6Ff6m52I75WRI3wonEIWdsRClrQ00g+GddGF0Ork9QR0nT2HQxquhL1Sr22SGmmNyBTS0JUu+RHfIoSaGOPoV/gK7IQglnsTLeCLyImLgzrQ0xVwVmoZbwd7NzTG3ySPyNGNBYFc8CbEVlE+Pvw2MLHkdoRtF0EzbEPU8zMmuxNNsJFexZilDazQIt5LGmUKShTg5vRgxkpCg+jtaGzIVZv2JtmYyxdwXZ/fIY5fkrbyVBqsO1SGmXBogT8hiU1hB/r2PQ/PFJsJ8iD+w2WOhtRtGQwh1oSs5+B6y+7GrwhYDlMp5KSM1j9cmyJuU0M0N5MXQg0PIyac+x5aEveSejoOk/ImPYmgauUwTHNGl+5jLZ/nFNybMGjFCoWRkFBZDw8DXXFFSGYPDG6PAl2xsaXRT3wUb8ASM/wBLJR6CQqEN7LJ7FERUSXIl2a/BB1M2dDCcg33MYNk1oZqSGtJ0GFyWkujpGRY0WqJk2JdHeRBro39j/kaXwKcNmF+54lkSroZJfseM/kb1OpMXmiUmfwZTXgTTw+hNVGSQSl/cc8iGtC+Rd+CooxyrRF4NwsQ2YLg8BZiyHkI7mE2GfgFBw/ngbpiD9k3RWQcoYzXB19hPyY00OscjZIaY20YdmCtEhqW3YY9vDI2Cduh6hs56IHl14GRceist/IYDSjfyhyiNFmyizK+jwSlNSy6WObSo1WGUUaaM0FmktjlsaKd+RuCeC5Zs3StGXDPjJUpghq/JEoka2WdFcGSuza0PYsIpi0qX8lHBghdTyPvTtkQivRtHoWh06PI+6Y+VyZ09ARWC+tCeBPOR4ZhGzyPWxdCo3+RjeCqNCwhuq0TyXIyejQ65/ZDCf6WOilFrgsRP3x08Da8mpkuJSihz0IrnZVL7GFRmi9ipDX5CIdtFDI9BrAmHz7PgVt5ZXDwqE8HyHrnQTyo8ju1iteV8CH8iSlpFJ+AtQS+C8oTb0VMvQmGipE5vgksY1HFEi0v5XCiDLY04aDePIth5GPD5Cw2UwxaMtMj2H7GP0Ixiigm0fkQo+Y6pjwWlh32EqBeYKxZJ6GYh9jIiJ+xvBT6IeSQmpv5D/hAq+Jj0WuGldQfKXhDpdIsOo3XwebEt+TPsn6Yg5bHhvZBg7WzB8DEsjcfKDrH2uPN6Gu0xug309I8BRm0ukNz5RsNgfQ3z+Bw1wZ0YThIsKirfRnyOjCZsYsup2JmfY3yeQoWjnYmSnRgJUzNGIi7RhlFg/gzy0dZE0P1wYjpQwDu0ytoeEnCixg3g9uMhOFKUjb0F/wBTuQnKQlwl6JkkErO+B4R2khu2LVIbqFAqZgVIXViaifYateRYK6K2E0E3h+B/gQZ6ExrRO0yLjeBMGz0aJUgdyXyM0PthZaRLM8iMY4H3OFGEP7BfFwyNPJoZaP34ZDkYc8cmXHUH0EIsYaDEB/iJiY37gin4j7UH+06jywlBljyVgKTJZdBvNGN70PPKyMDOZ+wqs6EGj0NsrTYsZPDaZnAGQM8piJ3NvIk2e/4GOlXos09HZiN0/IjTBtpdFl4+ehiS6S7EdK5pkQ+pjoWXdWBzec8ODdX7GoTykUB3ZGda6Q9mQ71PZ6jWirwehMibyPPJ+I2TUhmUaHwGqNQ8FZYMPNsqYfIoY1wbCoWHkvBkJkXShBZCdtGU10PJGRnbo7BBIhm2MrZ6H9D5ZfRePJ6H+k8+Eq+MMyIXJ9gtoQYPQ8xM8wps6R5dl+OJhULYwMjNlxMwaY6F4GGf2Lh1Uc6iCmYqU3oJuxfsbEzxsDpIh0LL9iHmpCpl5H5WaNcfOyI7gULYys4MnlwrEL7TZtpfydDF9NAqPUuBvh4HRKP2HgfMSeui15KW74NvCKOsswF/sJFXZDb0JG5n9h/7QoEXOxSErTDlixMsH+RQ6HQ02/RCTbJXSsu8riTafEaGNbRUjyQxYaVp+hqBMf8Ag9R4EPZkaVGQNZ2j8jwNu90iKc9izDeKsXcKbCYq6ulGep+5lDuwthFFoTSmVHIJKytr2IQMx2uhO/IsjmHwjHRMVGGOiFk2tm8HgI4tmCHhosE8GGSzglGWl9lhBp6E6LuzS6FegeiUa0NeH2Ml4Fg0QdD9cvj1xjnYyn7AL/qd+CEpIuOhYINOkmRPFMeQJjYnBW+EXoX5GwKl4ExeBmvRgeA82iLwQzA4dsyWCsfyJGxN40X0egsKeRPdEp1Cl7HaSdwy55Y1CFG/JgLk9kZ70eex8QhorYsMi6nqO2M8fwQ1BpukzYzXghP+xDz2IJsDtipzwecThkKNMs8LMNvIlLs/N5N4NEby3hoX/wAGL5Dlm40SLkEq5bZU5VGMh3Poa1pAiP4FwaE7q9m0ElVZ7FWc5ekN/CjmmGY6P8CIN+6O0RB+ayNG2N5wYd/A1mifY6C9DklsWCS2mIVF5bDUtl3WNsy9jm00A0MOl5jOqa7O8MdmBqpdbHmL4giFGumhhtN/sfAtqNjSpYh0tHeeDDsPAnUWXsbFsbho1w/cbZSicNhQfIErSY2FNDsVQedDHkODsfOvr/YD/Zu5oQWeRpvEMCa8Ga/vxZaZMhB0hC0WJC0LyQ8iNKLJoSZNMeAyOxOPYqX2NMNiGRXs8eIs1KvY34PJDAQ92KGPA1ZQlcD7CcdCROkdhiFXehuDZIo75JwaQY08FxRI/A3gt/wejYmk2Kn8Hsv2Mhk8ziHX5GJCaHRNpO7EtISvYsTA2RGBnUEdma3TOZIzY9ou/I6ZZkdGetGAbNXDoRIWbCZvmfRgqkApYkl1Rsp4vY6pMvfkYq30HUiTjMMPqh0benwF94uDVjZc9/I14cRkHHSD88Vv4G66oq7HgVeTQf7mRqTD7noZWksltOV5G3k8gl2CaLZ90LGbVqldFop4iYNOS08EgjxW79xa0ZG19P8AAiNp5z2Fq0zb7gyYl0LW6MtQzG4vY32Nm3xDA1PgaNsjI2O8no9Ea6L53xsOUaPXHDksvInD/gcpFfbFydk/A0aE/R/AB3+puPIyQ5b4EQbSQwGgbZs2diWWLYsNnfC1xeExb8m2SNKsoaeLxZxtwYENDxHYJReg5J4DvjYie115Ol+CISd9IaKw9Dwp1YnSL4MM7YWVplwvQbSfA2Jet0eYTTNZ8kDoLGciUgjpYRgvQ9BVGb7HWtYNobXskbg1svkQOs9GAzWekJNH5ZNNtlGb9jko8j+3kx1+xVqmQe4ykzTA4+WOexTXhiy7NMbMu8lZke7l+xgXyJk1emSbKPeEJc3RiI1oOTm32bn702Kc6KzhN4wHP3mknRSDtmJ+xlZqfYyNPsfuNzQyf+TCe8F6D9x+X3K6/Yly9DXKGi2zDGYaH7cG42fcWI2SSoc7SFox7TIPRqYq00Zq2u3QmqJHvCUkMoGe7n/gmjkyq/sLcVnoNDy6HQ9mBRwuGJn3GLZ3RvITXyTGDss7GELRtFKWBFmLPGCWuxvkJeWyRCcPfD2PlH9kf6R3HsTiwNRKcWG/yNE26LhDdIYBqmR7LBGxVss6MuEGhi0PLtOjb0LBcHJJ0EWwP0MNm2EN6g/eJKNuYELBPGtmY7nGsIJps/yATsHls86XgUH9I3/rA41aX2S6Gqy0ay5jyRlEHllTA71+C0uxQKjzRlQlt8QvqdUlHa2OV+A+wZZdLoWGV8jRMjrJp7M2EdtViT2zwqJ6FWYYYolfyZoYfrwLQ2myt94Qqn34Gj0YMx9+xsr4G79mo6MH/Y/cTsbj1G8m9nV7My6J7GaQ/wBxdkvofVyTyIpF6BZeKOHK/AtUsEPG/wBxm2s6HDbbn2EbtPH7nnZPI2dOyZ5bExhsd4rLdjKOnoqexxsN46Fg0M1ejL7hfYh3kad7g2VE2+xsTNUxrjGSeROU2VNBBi0PGowaBvHhiF1k3gZxd3e50K29eRL/AAJv0YGhrB+xvZqHlwgzoZYJ+GBHsMS4MLixeUWllKXI/sEEyYykb4U2dcTPLX0M/sj/AGnmdDdCUI0xitLJlPgWmtnQM6XguToWcDWReiEHnQlH9Yg8MGBvKEzJteehdSpGnhjaS0ttt4S4UqTbY4OTJgYUYNfI3QOS4FgdjN5lFt8ilqqHj7X0PO976uMBSm1p7OjCxrHeO/ZQIzTzGQUcrY6ClFKuQT/FHhqMsH7BKtQicRYwUPGFcv8A6DHUHYqen4Zcc+SOTwZltqsJPKeyiINQtNwLEfuJpFE8oYNyeo+zOpEZEtsb0YpMlNnS2Vn7mIuD7RrobQxNszXsQ1nA8q4jTyYVn4CZPLwQhLI7S8fY7mvCn7rLjhBqqp9hNEvwM1haMt6HrYnFvYyYexrfkTdFZYXtDDdrDMt/3Fl9iK6yIyu/B5cLkZbE+UwjIrweR0busGcmXpjhCzpFT6htbMtfcWXgb8j6tDwj7G/8D9DfYxt3ZtnZcDAUNEfAjcVF7zGH/wBC51iWO6Mk6sdPPcHYWKdj1EQm1CAdORIZaydezoUbG2zQ4/wZIeuGJFmB0sGPR4zsoxlKSo7KNnwU3xKYQyJPofH7Ef7Tz48NcH3LHkyWRpgzYRcCdGShZwNnArCex1mpozLZF9qoJi2bOj8FTTHnoVU8m2JnKXgTJ1aWx9z70UYLla82NvsTT8goIouVIlPJljT+RdxD0Sys5EWw2U3V/gOxMh39DGhtttvedTob4JyNHV+xksHIjpDZsPoHUqZjZ47u7/AizWbd6I1kYq9kXssxVkp2qZ3fUIJ89iUiyZvK6JNra8IZZ/uJM2A07/cqhvoHpaabyFMTJzSGnE96UvwfLWGyanjD5L+R6fQ2hn2e1FCq/ci42eV8d/u8Dqt4Y2H7uizsl4Fyj9x3aZWqZJ+RbglYu4dwwfRhhnGxoauTLyKxxPv7HSsFreTPkzZ79CKtPQ8tleKP1jI7E3Hsyw8mTMHSDN33pGrfgattvyYmLTofwNpzI2hlDTbUZWQCbw2R5ejR15Y9WYNC+w1js0fY34D8kp/BbwY2UkkUZAi7XaGflR/Dsdv2IhAnRhF4W1mZeCFPzZLymkoL7onTQ1PATjwO/ASX0IUeSY3waiIPENlGPB7IPYzo0izhsfFKLM2HRl8OGxk4j7A/3nmPH0Lwo8sb0ZKzBidGLKyYODTowatPZ2IrtwHC/uKbOSZUYvXgw8F9h7FqcVI7t+SAbbB5pKIqDwhD/CL2E2aU8TCCfg7tG+CpzImeT6iKKSlZYmuHB2mt14I7W9PozIytvJBa1lFlS9U+5bUjXs+hOL4lpn7CkxTM8BmuZ7V7Jp3KE83mEWzzkJr4DLGbTQ0bz+40Mt+AiK7w0/sEM1ZJP/2Q27ddkMv2G3sM6YD70rakOgyfn2RSSy+x70yyv7jrD7FnkKtl66Mmk9BPdKm3cCm/kW10Pa/seDIyRSEwr90Rkb5jum9vI4EzMqKZuroao1K/gdpPSeKYhgsDrfnK4s0y28HZUfTuH7KqKW+Bkl4Ub33c5NTOjpx7Z4MPY35WvsII4uhKnsb95KbNzJJV5+RUwyz3ROukVPGxW6xNGgjweLZsasmRPLG4Ga3oxcG3BZNdjwrFTJDLZmBa2s5Q0Mmsn8/yVlInmvI8lBioeX4FJBRqqXFekMJ/u6HaSs7HL/CF+C7koh8D+wxPoTah3o/JHeBzhi4OzIjbGLJoRrZeeil4vFFH0N8M/BD/AEnmJiKznoWUdFLwnkyoJ9MT6E4xBM3gjM2VQOl8gnofYesGYqzYMFaJRTZZsmAmsKwuDU9DeOVD8iyhUoFFscNmpG9s3NyEHr4ldB6EtRQ60x5uzxo7hr5KMi8Ui9/ZjaP8iddCizbGYHN8krmCB/LjQL7uGRADm3RlfXyQSnZgoWkWBKWQzzyzCEpfvlCQvDy2ORxl3tFqktGp6XOxk3glmtNo09nyyPlWZnk/8B/9UYETBV5Z4KRUm9Cc69i/cVhIQaGU1B9wG+hUrrEn0l7GsZp3FkXpDtCyRjpMVu5+GNE/YVJlNBjNZ8FU6Wzojuhpf5Mb00spBvXYkOvcHh3aNx4Gg8aG7lYYs4ekRSRdsUTO4LyZm6toooFv2Jl5/JpD8nT5cKbxg0qJUXJCKKl8mWYb1nyYq7O8iGtC+wZeoJ5Gssj8D2fIVY4jUyMSBuLSeHBEyqWQXyI9k0229Nicyx4xLHDy2UQZpCEjpkC1jX7iX4JEWz5kaUvsbgNKbWxDw9C9HV0KieR4PuNQ74yidy0PD8obox6hYbLOO+No0dFO+KUuC/R+yH+k8yCxkcuEPjYuE4ZMfpm2JmQQHRNhMUzmmOsvHBpfA3f8GBQc1SrwhuiqOjdwfxOxP9op/PbGV8r2P3A3WvCHHDxGY9DRNEsUNhRS4FKt8PA14GpoRVEN2HQW+GUabw7MXkdjW1UWbT0ZtyOvimw8ct9jJsc3lortBWCzLqgvulIdHZdsqkE9G7UYqYT8s3fVKSbO9wXHgbTSo7G3ZkjJWWaUmRh6XCFZza6S7HnFe3dGBwngsDwGZ2NNnciSwhBI2ztjXobEqaIE3ivRbK0IrxqvMEfwZGRjvtFFLjEyhQRafuFJor8lE1RJrc9FlT8QmVWQlna8UUurNDbd7x0eEl1BYimeh0dT4LdmStZlKLkqFHN+MMUtm9vyNTLwOiqPfkTi1gw+2LDjwiuAxpJC+4tIVvso8dizgVIjA35E29C5LnhkcwPT8CZN0rtE1cA0mCwxo35rt0G1hbbYuG9HryRXGuiSvsHYR4xaJ8ogplZvpoyC9RKVQJUJesDSGLeTLD0LTiHj6FxxeZkY+admnzT4KUXH7Af6TzF9pFPZi/I+IO08luEvSFkwNBCE8HQWwnroeWyuGl/YhNCLA8PgUkQdaNFexs1jMNKKJCGYNf7mmQYabznwNhMUMTC3sMZ9CcYSNaFpMjZryVYf3FyoVvInqpRRHTtBMknhWvBRLatfl+hndMeBQkfhw4N4FCreRirFYf7BWuT2N9kttiuzs1k7XpH5adW2X3PZUMbYiST7JeBVG6v4HkbjY9Sgsz4HrayumTXOE8eRph7wiJoTd3UPJx39zWm2IVBw1tkvnJsyqCGyvSG7Uv7knGrsTFt2GRaeDd5Yoyza+dGEHsSU274En8gmswvQtwmrn2HhmydVuMtlYBR1GsUrPJ4GqJl4Qoxc/Jh4+S4GPTYder7G3SLsE/CO/oh74Tq7hrDyOL2zLZDxk/1RdTaNlfJljcMb4sXsTrNdjysFeAm1ob/iFDqeMti/zqMpSjtkP57EJI6vY6dQzLwWaJNsjdXMfyRKxaaf7l9pyKRGSfsXeWKqVjYmd537G1dpDIQvsbGytaHaQVpsYpObw+Y048PijJj6KLhn9gP/AKncac02YYsc0XC2Ubg3BMja+Rs+BPOT7iHl5XgSJ5WC6fsYHmkrLO7EJPdKj79wnJ4MM3VUg5njyb9P2aPdHW2K9owpnhG1iIYsaOraIfSY88r7EGk69setMJ/Yu0VHmbemZKnnwZSYMt+R3UnTwKLIUs9WWeR6+vQrer5MgSTMAnrp9mytYY9mtjz6RR2FwwO56HtnJh2PQbE7UbeBWsTwywqNLBUtvxSRhGsO3YpHOvRX5mkZe5KR4jy159IyFX7TZgTJZWPZJJqVEaa6aRhCsjnui2knFjZlKmZmklj8BtzOU3kz8EynDCNrP3OpG7M7abeZcDV8vUN1CbReyRrShdiBV+RNYf8AJZ1jt0bqaIPG+/AoiqDh7tM1FnscxmiHwPCc76MX0x4M4suyqkmYNpfllp2TNyQu8lVMvsXG4hu6wOexj51T9xxwnjQwneFLGfMNryeKcNrBOsBGyteP96HNVVSuhiMnbfsXDBJvsz+wiWddsdCCo+mTXQumlB+xCicG4YLFOI0soa2PkWv0KaRLX7jS7NGTA2YI2RCRqjwZG7w+GMhM8XjRv6Fxo/ZDH/czNRwnxsbNj2eiYOvpbR1wsjmBSscMoPbfY9L8l0Lc9ku+jqim88VZUbSmcxdyi7Fl6I7NWNVe3oTZQ3ik0xVnilN0zW4XgXT3uUFmljdvYgLizXWCSZu1DJHVLgTIXYoJ+sJlI08p4PA8/IjL1Z9xjV0g6aMbMJ/YWEQkXXZkwJutHQnlk1bI1VDpOVSK30ZRF4G5x4Ji962YMQUmrSWhS5XmQZ01fyNSdcdGsBG/FGrp0PdKw3E8FGG94GS3EVFO1eddEF86RbM7ZqZEkUj7xgwiM2Yo9CDbnNKTNEfY0o8PyYwJnpjVfIW8foVZPo28+BFj2Kbwiq+RSU58dnfsdVu8kIl4NFOxvgHkWFzQ6bo2z5DjgVpseWPGdFfwbGrhMErMWoh7ZjwN9jeA7hs8hABdv3oVqIqibCUH3a/sIJO2SuzS35G9xv8AuEgybuNyoRbRCTfoStwu3YwD5fAd0S2mNT2hKwaqCUTGRdHYmqIt5yN14FgV4DeDt8b+hjEPhicHs75Tg34R/9oADAMBAAIAAwAAABBZWJzA0cjPSQZtE339kkkkkkkkkkkkkkkkkkkkkkkkkkk39mhF2AFNt51mW22Dt0wWB3nCgZDbI9/t02EA2vm9+k+4J5QqCFkahH/NkKd3lkkkkkkkkkkkkkkkkkkkkkkkkkkl+30pPBG0TRgamhko2mlGhSD3AjQARdWdfvkr1Clsn/l4ujHJGi1k3RXtLGRDq/lkkkkkkkkkkkkkkkkkkkkkkkkkkl/jwI9r+ALxw3u/Mk008vG8SzLvRQQbUrZt+pKgr9p9fiv9ypb3Z7AjL3JlCu28kkkkkkkkkkkkkkkkkkkkkkkkkkk30kj2t/MQQLq2O5CvGmk3RpGkiMcCGNUYTLUG/sTvcLb5xcwIoBe0Im9LfLgu+/skkkkkkkkkkkkkkkkkkkkkkkkkt/gQBkblfaOTUj1uo0203t2u82UF1Spanr7/ACQWT72U7mA8dAuHEfvOlp4mYj/97JJJJJJJJJJJJJJJJJJJJJJJJJJZ/LI76wSBUL1ZIrbW7pP5JNorykFGBgJG71Y8EG77dD20QNJgSoSfgz52QYMU8/JJJJJJJJJJJJJJJJJJJJJJJJJJb99CxEi0GHQVYfX/AGyK6be1smSwsrANnYVud5BpohsIM9MIB3JuQD31tmVSqUCrf6ySSSSSSSSSSSSSSSSSSSSSSSS/6fEM9lIJNIK06H+369k/398+TXs6aya16skBtBksMFJJFFg1Zn5IaBf0ikk4txeWSSSSSSSSSSSSSSSSSSSSSSSSXfR2MXQlhslpTnYA9m26G3+/mnjHFjSaamnpZwqNpkFFpPe6bVjNJwACTbJIUAC7+ySSSSSSSSSSSSSSSSSSSSSSSS37OBiCF4T2lFX3A21n3Vnsu+33lJaksSbTQdfYLhBvF/8A72g2dq6yVffP+wSHKNK3tkkkkkkkkkkkkkkkkkkkkkkkk/1tDTr20OpYdvmNxfZbkpDLTZ/9/vKckW0u3iZYG0EhliiFBFdFqoG9mxYd13lNv/0kkkkkkkkkkkkkkkkkkkkkkk/+loYHJP8ArbEVpf0Jl3z/ACxH1n3+2++hIlTXf7wN/aZ//wANiiCkvvRZIz7VmJxU4fm8skkkkkkkkkkkkkkkkkkkkkkt+0kDUOJ03uzTmtkHAB79Q95S41m89/8Afw265dNLNLbZ54u4VMsp58XAE4AqMEXOff8A6SSSSSSSSSSSSSSSSSSSSSSaf9SFA9sUD+6ENS5qiJMmjT2//XaT2SX/ANmU0iDOa2GRtynGM1M6reN7LbwUMBAKAX3tkkkkkkkkkkkkkkkkkkkkkkk/ztBl6D0qrTJcvEMCXprNQXv+39vn2ns092pxFdkMWYLj+Vos+2msezWAAC4RJTD+8kkkkkkkkkkkkkkkkkkkkkkkv9/LF1of4XtjEs5rVjyTtZ/yv1vs1vmmiwnKu+nnz902ca4/NOw0so5Z+QYe02uIf++skkkkkkkkkkkkkkkkkkkkl3+n3KFkF+iAuQknYJCCAAYLrG01t8nrMRZTJZaTeCPgLZf11T0qYtDHKQT8/oDoCE3+/kkkkkkkkkkkkkkkkkkkkl0/12pS9wG0CliSY5bKTQZQYZOYsmOBqBPFJcvuY2s+pKZsKorOk2vfFhaGpY24CxKc3/8ApJJJJJJJJJJJJJJJJJJJdvvl4SmUvjfeyirjyCmkAwUWyy6Iiyi3gEWXfmE11otuykEGZTtlNdbDRBPdtQH+VIR795rJJJJJJJJJJJJJJJJJJNftlrUAO3eSrJC2hTlUgQwyEgWy2mbFHKrk/wCuzQvpxJAFLCarlASS7/MFD/ZdAmRDzv77eSySSSSSSSSSSSSSSSSST7eaVtA+QjylXYpFP8tAvlMIFlt05v62eIkOTLJBIAFBFM1QCUBSTe+z/VEIqSsfZAyE/wD32kkkkkkkkkkkkkkkkkl+/wD/AK5BXdL3Uj6gFP3usN+7sskktthNyokYMsKolgJllrxvffLdCQXe3X0sBETvu/DZtneL+2SSSSSSSSSSSSSSSW37WvYRiRmHRQAXUzjDP7nu3hhElsIbVJa/cpV3kozJHEJlJHPCCwRNX7S6R+7leAm0ujqrTLeaySSSSSSSSSSSSW6fbH6GttmLf7mSokx2EUMv0tlkslkG+kNoaaX8vn9/bVBcEJ3lB1wYU4tB9btY6gfj3L4yZYa5byeSSSSSSSSSSS67bY7xQdk0XvFqC9ix2kCk1QcBFs21s98hv4YzaW+ll2vo40BbRedWJDkSbpvcHuor9YIJk/s292/766ySSSSSSSyz7/H6XMS3MO4vbjeBtBfxl3rdVIkAsYBezyR2Y2fksNCTIppG8c9HD+tGzTGzX3S5GzQT9bEH9MnL3rfeWySSS2T3/wC2e2tzCHnAVdJ895hST4/ASbQ5ZTUpT8YkG42uuk7vXbPsqEmzTJ5W09ks3k3l2t0JpLfvpHTfjLT1/W/u09ml9n/+7/8Arei1Jwh8OXMahnMRExkEkbXiGW14tMIvLcYyuB0DRpcqOcKK5Ci/pNbJnJ7eJHk7w6rCLQp5wm5v/wD/AOkt3/8A/vsDss0aSAZuMoW00q5ZYfnXatIeAgf7EGjEk+kntGAjKGEjZDPyaLbp5pB67N/bwQzIxRKICilTmCuNv/lv/wD/AP2y0M95QEl052ktfbSgfV2Se1OHE41fJqn0rlWOAtwrK/ArCW6E9b2mTMNNOk1n98jdkOzjSB78XbI9yOJu/wDvaoLOQokmAAmJLQgMB9+amiWmI1tVDJLdMevekQwxMxoOegG0VH+xoPJBLcswE8env3BJq+sHd4alf9kSues2Y/bIWxWk9hxrBq2y3exnNN5HrWyZ6pqRPNpqaQeNUXJccbxsxhU2lFnP7NIWk4OnfJ2+Z7ZZNYlDgHOqcAHtuMpwJtyzqQ/pz4lbUpFGyXEAjhpr1ea20qAvohflQcWWWXcArTe7fS5GpOOy7AIRZfD3hYAqj5O5g1KD6a+kpoN0cbtqQcwd5+U332Jq2cpipyIz6RhNIEPMKPCFrtbtk1tC+xUcVapxrK3b+Xp0cWRfL0hhfGU2iieBOrFEuKpl2RQRRpEfjXPlemX406xe6Eqr9bUvtW9gREqvjNR+mRNKjoh/hr4wMUlXoaLKI3w3WiCykkIwcFoBDADXVfuMTfrZ74CpYUtXse+E9wFLlMD0GAnlmduB77bbyEvU26pQnkMb1ZTYN9UkcSCh/F4oq5yNOv6dSbqz77i2zhKW7MZwOclhFWawN1bZrXaNjXb8dvOLQL2/wh+iXz7a+o1wkm9Ga5tIdqz2jfZucIq/RcxZak+EcdtvWCdDSCpGl+DFAmbL1sFoW6CbSRcBNflztXAPVOpIg16NBCczHyDLBrmEcF9ldKprVgZXIONUp2ZKF7w9ik6jZbsoOYfxI/IXinJLKYAoAEZH5rbebGPpqNech4y7duHwGgONS1LkDlGSK0DWQBg63KP8Oat+hauXPa4Zksi8c2ZIuYa6R1C6U+AIF4y0DM1sjKhv78dZSy3VtdMdWoZxPUAznel09IlsAEwm622qaabyuhCKxTqubHm46HZnQ1P8do+2oLTRwx0LI3CVWAQoTPwQ1le/rQqqr3NnPdlXnc5YXPk3FYndP53ZJi56WkZoiQe0UyheDUIoJQlbPRnhGYbOjGJHJDAiT6u932USveD8OXC0zx9a/YdMfrvIordvkN3dfXZmNjnd50+TqiDwzxPlsihMKYylVJQsBw5pdXfmD5fOniUYULdfFZxxEEdFBGMY1F7RYtWiiCBeGRTn/wAJVKba7xNT0/CUB9YK6Fot5en95AIwLUuMGbuu9GT60fMPvyy2Gbwcai6U0WV/hmx/RpCANCAuUK9FNRs9FSDDo05esmGeIsfSk5WCddjqGTVUNdm7r+3ppbVU8i55JjNFOBqZjG2SeToHHiCR99Bjqz/jXN6TlvourBGa9VAk20xfZDEviMYA0FCapXeC3qQBuaYOEbxa2Rncy9yzW8bhXl0g6lmiiOYqezx/lCB/nY6sBXnf33OXFe9XHA7ghOSVXg/kqh9VBIVH43T82HP5Oc9v2sUb4Fnjup1yxnYC+dOWxX5Vrm+YLR3udJPow2BYvX+Y/MW0QLoZd/Xjs17pF23z34mrwYuM9JIsBMhOYzvq+Z6wFhz0obPHZ8qTkDj/AOQE23pFRE1JCb3GhDqEkRaH6VQT7AsuX4G/YX6M8vhsfDhOxGj9nAl84FopnqFP30K5mNHDpvghNA3NYxGU4nJmYOBe9vShWRxh98WRPrM99zrnZCJ5Kd4ekF3kusSmBOxQM+Ir+FzdHAlcZAvNH6eieB91E7PV7OIsDmw10c7/ADbGd7pEopU09WoCp7+Cj38Q50Wz5U3C0EWhUCOA65g4JsbEUTJGUXmzR/6v6sxi5aH2YuqW2xznGzkgSrNLC+CFbWrryui5yJQm+KbXUPvOmmbVMVcoTD0U8ROutrgkjBhdVmSIUfJ+uBXuWe7SzKRnYBYvTIOpWHSkYYjyeTga8oV4P2NORb0QN8wcAZhl90S4BiKEQS0fJeMm3tlt9nWZOSo/HUyQarhOhgwG1V11wzJrSCbeNI2nrJaccGJIKuYc7HvZEHiiB4z2dTloYKX4nz24M6ZY+4c35P3TlPHShOndqvlF8psrD2kT53qBL7WLfdqCl78sHHkgafHU8ydybXcu6otAiZuKFHyhtnhYhIdCVICFtS35Xfhkhv8ADxSyp8k47v6wkJlLE+qbmc7v3kIXCIRUpCnrm5H0WTD/APgIcDyxH4tGxALwIj4f+1pdbIzgHIMSfxhGmKN9D+gnWKUh+YHKTHCdZiGCYDdl6t4puaNBJWpD4ngUHiOYa3poh+xeTad5/dZNQg2hSxgHbtQAOL5gI8xUk6PCHKr2YA1uQdd1Q2X6qpPjrqpvpeoO1ww6I23AyCSgFHdBgwzVpK5xArvF8cH278T1Vo2KEXGBBbRbcpAPUA67SYNIbjfvxIq0ULp/cDsqYEwErDKJGeIEoT5jlbsYfnnhWuKSPu6PgCRYjaGmEwpwTxJD2B7i7wtrjxPCe3gcM/HkObWR7+kTWvpJ03CEg1XLYW/+y5qTSA+7HJtJBNHv7QWrAABwUBDjM3zW2GPWsPqjJx59pjZfwTo5kJVdGaSxS9543urZO2WBBUly1n7lHGTGL8as+ihe3lr/AF8m2o1gBQTrFTlWNYTCWCcOWdJp1NITig9YJO8KF43XSGX6eVfeZyfCuDrmMn83B6xwoWXRtU+agIEGT87DVokTzsM1oS6x0+3EyIMT6L4pfIpeQfPIpv5rZ3ckCyR37hf2IMZSxBikkN3Buq/2UTvUf7HueKkhbOQzyu8Li2Q/esa3xWpgRj8lKrW3TVus49bQnOCsTVN0LrPiEaLzq6TehAZs4aFRkcklC4PaSDwjT9cXH7jTxJiWdowrylatnsw9/ZUPIm+cBjSYpMtI4yd5+8sRfA+DUUwK9nx5p80UtcLlBr1pmjkJFioBEez8T/1IN5tueqoHnoCmG5OdnohBFpZJon6agZXJBCyedJejjP1W8Nymakui/g3OKPsLm00NUYcj/gwMib/DQtmDkOP6JpvGdTT/AAU2ZbviyIXhkBY5BH1JpnY3DYiG7ze5mwdgoxzwbjiETbuP6mBvcQQm8nzL2qsp/8QAJREAAwACAwADAAMBAQEBAAAAAAERECEgMUEwUWFAcaFQYIGR/9oACAEDAQE/EP8AJm/C8PDzRj4P/wAGsLisoWFlYX8J8Fxo/in85pn+TD5Pi8MYx8Hhvi//AAaFlYWUhImVwhPnnJl+XXxQf8Fs/wAmHxfJ5YxjHlj4v/vLCyliYhMpYSwuS+elL8E+LsnxXM18qwz/ACfE8NDwxjHwY+D/APBLCFhCwnlCE83hM3jPj3/Co+cIQmJjr5f/AIf5s3MOsvk0QaINDWIMhMT/AL6wuawuCFlcHy/r+KsL4ZwXxTlOf+bLwsvM4PDwx8GMb/8ABrisoWEiYhBcOycWL+Prj3xfyPE4o75f5PlY+LGMeWPi/wDwCJlCyhC+acH8L+Ff8Ccv8mHyfJrhBoaGszDy/wDurCyhZQiYQuC/gdk+BYXGYT/4kP8AIsThcvix4Y+DHljy8P8A7SwuKysoXBZeZ/FWJ88IPn3/AAWf5PkmGPDeWMeXxeH/ANpYXBCyhcF/FmZ8MIIcENG/jhCEw8zE4T4v8nCcWTg8TgxjQ8sY8zDX/ZXFZWVwWULjSkzfgnCZpfih6QXxvO/4P+b+C0QZCEwaGiEIND/8GnilE+KyvhfCc2hcZ8j/AJ0G0L/+XF/NMQeXh5eXh/8AcWFhCwhYRc0TLxReHRcMnKGyfw5/BfKFw0f5OT5vixjwxjGPLw8P/sLmvgWELMJymJi/8eEzPghEOkIQb/D/ACY7J8T5Qaw1hjHljHxf/VXwLCysrjRcaXhM3MJ/NmEXH5yhKScJh14fZ/m4P5mN5Yxsb4sb4v8A66ysrghcEL+NCfLPl85TivjZ/kJxo8P4WPL4seXh5f8A11lC5riuCyv+EvhnOGuC5PGhn+TD4rg+bQ8vDINZaJwmZ/1llCwuKysLiv4k+CmRevBR+F+hWNumUuzrC5dj4T74aL8bNn+TD5wWJmZaGTEJhjQ1mD4PL/6SWVlCysLEEsLiv5EIQbLeO4232L6Ho7EEvsbvwlifDCfFB9n+TD+OYZcPg8vDw+D/AOslwWVyWVhcrxT/AIvRYTjpohMEmxu9FE0uzREQhEaNFK+Mzr5nT/IsP5FweXl5eHhj4P8A6S4LgsLhcLC/4PRZhC7H9jc0jZSlLmsrKUpX/DmH2f5Fl/Ix8GPEGvhfB/8AVXCZWFhC+RYhOM+fouLNoahf+C+z/J/Eebhj4PLHl8H/AMuE4TMIQhMQhCExBIhMQhCEJmYmaX5uqmblah/BBfHL8SGLD7P8hCcF8Tw8v4GNYaxBrM4T/kTjMwSITEIQhMTKysJcULhf4XRy6Hb5ly6P5mz/ACcEuEzMwhMtEIQhCEIQhBohCEGiYhOE/wCJOEJiEIQmIJEJiZmEsrguC5VFPBV6TjS5uOsdOXRjdwviuKd4WejLymOs94Z/mReF+OEIQhCYQhCEINEINDQ0QhCYhOEJ/PnFZXJZXwLjS4peFzRq9YSuhtLS4xn6Il6Rvok74trl0fyUpS5onjox8KUebmkZ/kWJ/IY8TDyxomHhky0ThP5c5LiuKwhcV8NxcXmt6Eq+huaXLwTTVErg34h5Zf2U/T8j8CPKVMfxQSvQ012TO+HVje8UpSlzR/Y0NOkOnZ/kX8Z8GPk/gY/hn8efIsLguCwmUuKUpSlzSlKUpS5o1Y29FKUoneZKVfY/bP2EvwUXSL946KyijT7GuxDC0VTZ9R+Z2OcaUYW0LWkMMvp5q/WR942jQToNRx5gneYJds08G423p4cOhs/yfw6UuLhvD4PD4PD4Pg+M/i6LmEf0fgfkWYusZN8PQEjbZ+wvtG/rQvdiW6xX2X9lfZX2f2P7l/Z/Y/uX9l/Z+h9JDwfaRteFKXFKUpSlKUp1CYf3wJJdIpWXHp1wVuxdcJB43c6RGysYjeDOnuKRIUuXijKdjpRUKvobFePRoeyTC+sQ/wAy+CE+B4uaUpS4uLijZSl40eaXm/ljPyPxKYSvgn+CZ2z1BKCX4Ekus3g/47Tdobe0NfGPxI+DT4RO1mniYo9YleELov3x7yuL3WOz8PcTHedaxcvPuLhkKeYpBjw3hFxcLohTY0Nn+T5aUpS4o/hfBjXCZZCZfwwTukJoT/D7WL7hejEkS/BL8Ejwnzy4eHynzznRs8G/wXi+b7xWnn0TxvHZwpiXLuIh/mOj3MRcMvg+8PWEf2P8x4Qg9DTvR/mF8d5XhS5fwMeIymqkU9wTukNXaPyPyPyPyPaDb6GrwpeEZ0gZ7cEO2JYS+kLm8KUpS/I8L4JlfIhfNRCXlS494+lRT3FGIqsXfDrCWNDOyD1tDVOtC7EPRd4m8M7O+iXon2S7wuyHWGf5BfBeVKdAh/UabMBNNPaP0R/YaeD9D92MlDooIOiJ0iN2hJF0v/w14iou8UpSlKbNlZcMvxQhCLJCEf8ADubzXwJ/D0UmLnrMGQ7NHp3ll3iYo1j8N2wIu8vhB4k6Er2RntGMY8NHguz8FhD+hIaeLhob/wCIv3LHZfDIvs/sRP0i+yfYg1Fr0L6o/oR9FX0izwplKLzeUXEIdEuZyuZmYmIQg1B64ThCcIRYTJGT4e+K+e/GsvjLiQs0sz7wiCNHpoWym7HSc+zrDz7lkp0U/vG1hHuGtHlKIQyE9ErGG1/okJo6ysS57x6TlcJ8Fz2M3hqiOzrF8KXJ/QTKWFO8PPeGqSDRP4UIiMKKI+cxczF5LCEP4bl4bz3hnvGFHrhcdGe8VneG8U1wohuCR9HRI9oK1RqNfCqJC+kJ7pdGzKEzUb9hSW9G3CiRf6E9hocKk0Nbs0iJoWuyiZSsrxRPjCE2IvwPEw2uUvC6wtcEP4NYhOEwv4MxCCMlEJv45m8YP4pScZcQ6ZITexog0NCSEiNqQmxaEhtLCPoeujcUNn6Vp2icbY2loTMTOxj2LRKTfYyi2OIqIRBsNvGjdRnYd7EzaGtSg1DcSJexO7IQmISLCIJCWaTisd46GJcnxfFYg1zfKDOvgnJfD38OiGuU+KEzMLMHmEp0VMcRcGz6L9G2tjYM6NtHo2UipjSZ2oVC7G/II/oVdCNY72N0pSpFpZhsdlQ23norHoNvzGkNsEeYhD8ComNAkQ9JMT7ISEzfhbKdYTx1wY2Pg8LCXxzN4P5b8Kzc+8L8dxcLCGsMQlSE4axcdIhKSHg2LTGOhOIlEwtkG0ejiZUX6K2z8FFscR/R4XCKJfZ1oezd6HtpDgScNtjGqimKexX6SCltCCaUZqCpMWP6z+nuHhIJ3ZNjWP74TExM6zaUQbpMUvwTDEsTg8P5pwn8FYeLifHOEyhFw8MRIjoWW4IpDQ+yEo1MPGhpMeiumg+tFqEfoyDRKikK/BOFQsJuxv8AYknYqSItgiBq6ISBo9IojQaOiVsSpE9tCR9DvpgTPsb0PK4dEP8AeKII9KLR5s95MXDzFHnofB5f4ScpiZX1zmF8M4bz2TMx08NpKs/qLZCEKXF5IfLvCO8e5vDvLGIuEW4eExC4o8NGxLBe8X9hU3sa6ISp7Go4VHXhtnSEu0KIqDe7GkMcsbT1CRBprAyidkO2MSkJRux2ejVCh/ZBpEJdYLpHZ6NsQnBCzMddimizMFhFH9iw8TDe9DJhQexPk3jrFr4QnPsly/hnyaGEyzfOCGiE4wkeViCwoPKOsUexLGywZaam8PrHhREhENOikPsfg0cGqjsI4JXs8mNocuxbQohA1FpjXYtCpj2SItUIhPAxsVhs2Q/A39ipFg2UNqFRrsq9KJ6R0I/sjEhQSEiY6E0dqKNDQR2OWJWRlkHxQiEEJaNcGyjwnxSH8Szc74UuIT4lhcGPMx6e8PefeJjoeycEzsedHSKI3ho6wjzCcKmLQ4JDeFLB+Boxt0rbEUEfQmxNeje6h2WiElRykZ5BiqdY/saFoiZpndMRNDdZS1HhIN0poXRRaNMWuy+YWxFxGQ0cGqDQ39iey15aaHR6MYoWDezofeFs6LweHyuLzeIb4LE4zi8PKzCYeaPnrh2InBuZouGzdw9CwtDztYomNjZs8O+iCoxP6G8LhCXo1TQbwvTJ6xNdDogkKGN4X7IrRwgzpBPwsGzKLSOxVC17GrolYkwytnbErpEQulhEEPYhFL4dYYmN+Dfo3cEJD+FaOxdFG9Ggx2U1lEPRDmHlvKWFv4X/AAu8Qh1zQuFLi4eKXeGxDRFSna5Jcd4b4N5Z0qLQbUuNTeKJ3DwVdmizBfQmNpMbY0/BM94OjISFRPodSHDTobUcMY/RUxtjVHHoca0IhKBKoNLw+g/oXcLdCERHSELRGJaRIIRsUKLKNsLTz/QtIWyRCQghPQnjYlJBfYhivDrDw8dZuELXyQmPPlXJ4pc3Lw+PaNlp/Y3zuF+4vBjZ0PeWdj6NJY6GxXorR2UUbcw0MajUKxDYjemXcExk0I29DRtdC+hsbVLh62dhwzsekhCCno0vCfRIRBoS2L2RrQxttCS9IWxoJQp0VLoZ/eFRbE2jbWhMQrRMJC3sQpkEo1NFGL6RJ0MbuhCFRaysIfGDFrhrs7z3logsz+BPhnwzELcoZMf1lDFi8GVnQ2xfuL9DaguxFg6N5mDOkJtFV2el8NFII7RsILTHQn6VibNwSXo72NBxs6C2UuzskJdk0Lo9hGjvssZWJ+CJPY66IMSDYnNob3sqD62WbKhWIehC7o2IW+xpCX0LsgiKjHpjS8HOSQvssz0R2aMTnRUaJhaFtjXCCZTsQuijKLHTHBMZPTr41zWOyYYyYpc+nvGXvgxZnCGyC42DIQnG0bHGxOj0f2UaEx94czE0SHY3C7E9FwhQlY52sJDaeyD6NkIThN4aH0EyGkfTBQJNi2EoxPB7J9ERSjYn9FdFxp2MWje4Jr0pSSGqToSQkxKCrY0SEFoSQmhemOLUHiGvWKw9KUv0JwodYkI9G8OmOY9wnhYkGNZh0xiRs7EuUO80Y89n5icWWZWGhMuy4XH3LfC43wh1iUkGx9YeOtD0sJlEJlNi6I++EHo8wg+jvHSI2hHbC7LBC8ng3FS3YmUdhBuGhUhtibpBDVH0D1sT+8p7GxOvQxl1op0NsTnZXRtPoT1Do9HiCRsL7KJp6KJzFLo7EOhfaGkxNC00wTKh76Es9G+haFvsRfHiCwuUw8w7G5ickXg8K5WOi4WGh5XB3HWPS4gjvFhc6xCQ7I0LHh4bzCZabGUQiIlIxJtj7Hhsb8R/Z0MWj2MQaSi2GsXw6GKbDEM9K5sT9NOxNrYlTNx64u0J/YmXZQcDYetDpGx6UHfMN6hS+iYb1o/RfR+BNIoo2VfYloSh3hEEnhCJsRKNIb6HXZR+DQn9FhU+sJ+FOhtQWuhq9EhRD7LvHmFsgzvNw8p7PcNi4dcXi5Y+xl2PeEXDx1jsVGPguxnR2dF4LNKbYLBUdFRc9CWHo8GTdwqQQgkhPoag8XZaMuirFEdj0diGMYddYWmNjK2NwWyi0tdF9KxBPZazpjex9kvYkGhDtsfoR+YeFfRrH9YTLDbIdMLGjfSGRdn4LQtmiGOynsG50bCtDP0viEO3RuHZaK5ip1sv2XHmN5vmEKDwybIPEELheDwzvP8AZKx5os07wtYg98E/Bo1iYuhdFxsuHhCzvFyixlGylwvoKypjClEkhoaIqmuxjuNlgq8yos0eYTvZqjPCwsH9lnYtoe9rFFUdEZdPsQLfWI+xvw0cGM83hmx/omXwZVnsZYUTRQgtoah0amJWejRbFs7CY2Jsh0tCW8JaEJlZb0LZS0TKUiZsVKxbw2dYa+hcHjsmOjS4rD1in9EzSCGlcdkwn941hELkn8UmP6IRnQ1SCWFoeIQWFi8H+HQmxtiZBX2hWItfSLYh4J9HtoaUiMbbKmyJinRC6Pdn4M8xS4XY2fpse0KjeUXYnBIhLYShqmjtjGqOD+x7HSHWf074LpUgibp2SERKsJbo3exPUKmie48EJ1jPBfYt7GJbH2dItILs73hEp0TQsXDOsdj1h4mPcTgy4Z2eiE6dY7Ef0OjnR0Lj7MPgkL8JxWtmhBogifMj3l3h6wx0T8YmhDVGoegii7fZL2OTRD30JRDq2NjP7KLZpY0NDSTFPSPBn4P6Kusf3hCG2sNA0Ymi3aJsTZ0e7GRwixcdYej+jooTcQ3s22OKJmmdI0ZU0bRR9iF2dE3hD08IT3hEqz+cF6G9CKWFEX6Fx67x1ibOhTE4vEx2IuGO+FOyDRDsf4bxBkJlEmPctm2IpS3CISZXxvFpaPYod6GiHRT0/BaH9hSEeh6WjamJGhq9jWhNi0hv0bo34PFmHtnQ8U/RvUQhpTRNm4dY7E6inh0hMUxiVj2QgxpkNCbHp4fY8w0I9E4tDdEmbD0OdnlLR7IPTHWbRtM6Ed7Kyspl2JwTaLRfZbjseiiGhLwc8O9CLhQjfR/Zr0vX1ieiTFrj1ifI8o7IUnCcXnsg/wAKQpRZ6O8PMEsbzaTL2Q2LC1j+j+8MbLR7E32J6JNHibYNjYY1RqDWqQ9Pw2MWWUWisQyUa8NLHR2WCei7EdCcK06OtCQbvRTvaxomyD0Q/B4rF1rDeCUI09if0Wd4X0LqE+x9HuKnhCX2fiEi1GJwbghaUctDtCMmFsagmNnSNs7DQkvCDQi+nZrpEb6NEO+8dCx3h57w/wAOycFvvhCcZvg8zCwzrD2WZWi8u1icLXlvXDwuKd5bpPMV4uyicGJbI3tFvbEwb0RiaVjxHobvRNVi0Jzs6Y2UeHCDfhsrWhuj0f8A3DY9iwlVisbEr0JtGmNQlKkhpM0z2P7xBdY0toSYrTNlBmWbH2L6Loo9mph/gt6Z+C7VE4jNGdmk4yV032LsjusrrQ2+il0J7ExUNNCYmmUb8EiiaKyJOlPOEuHjWHMQlxDrEhMwhMrMLlMvBi3nWUIZMT0ZZi+4eP07RuEpvCGWjOzpYRT9JjzExTrMR9g4KNjVBJ0fkT0a8JOjsdQg19DfoxI9HoQ0lst7KOnWsQfY2zyliKVDY9iZYNi2wbI2dkUY1ehkPzC6Q198FHBoN0b6pbtjcKUXQvpkY3sTuxK9Fcg9sYVdnqg9aNNpo6Y2f2JtLQ2+zsZIIuyjcExdYVP3hfo8ymLeZs/CjQhrD4dEPwTNHfH++Ho3vPZCZ7xCPCUz3y/C+YsNPEG3hMbo9aNC0dj0N4aEdHXZ/XCibTqxSH/Y1lQrbor2GW8I6pQmuy/QyDUwnGN7KaHMNwtFo3g6LZtbO2y4ei6LSl9LiiC0J6HoeHh0E0kJJ0W0eFbE8Juiot9n4WbExOsmHoNhdaEfonVsSh+Y6ejw0LZTp7NBOouC+yluF9FuhKI8xS027GPesrWKUpUd4WFs0svQj07xTR2P8w8Qnoh4SxCix6d4uOi5WUMaEMpcNvwb0LHQ94SOtFQns7ZdjQ/rDvmXjY2yHmjf2PKY0bY+iEsjOxYzbfQ9Noe52kJHpiNdMSfon4PWsaO2T6LC72ddDbeHpaK0djcWjrD0dokz7iiZS6z2xnQgvs0n0PCdYvobFUKUa+h7E8E1VjdG7sWhuPQ9liRth/eLgmkVFG0dj0hF8NNGw2P8FhN0p2P8zUdnWGeCdPTWO8seKN4n2VMokQqzTo77xIMgriYmaPFws3Hgn9idN3L/ADCeE9Gi/Y39FKWdZah6aHsZdF9GUbIUr7Hi4R2RF8G7M2dIjB3pMToIZ14Im4xKG/8A5kl9kbGbHo7HcKpi3WNDWxjw6J5ZS/YvzFEemxNCdYuHA8aOjXYnSwWmEWdcD2zeF+DX0bpd4V9F+i7o1UTGx/hGuxha1xWKUTojzRfvC7LllGd9Gzw3n+uDx2LXCEIQo8w90N4hcXwSg8zCx0IY39HaJM+CYyzHeFhbJjsng9Z2bY3CIRYtnZpD30JuFHiuo1hSYjXsbVL1ofYbMdbgwb9oSYxND0hj+itDpBN3BorGsMtKM6ETcNFgxLC1ioWKE9DTZ+i+ht9o72aF+j0LC1hSlEy4ThKNDpiYnsTSG69nQ0EE4ypYMKuxvo4VsbpV4dGxaLBNFvZYO9lKd7Gx6GxicEy07KI0Mf7hlzcUbuP07y8OiYy6Kn0QhBPHZMXi4aEPssEy/QyU9EMv2do/BaZasLQ8XZ2zo3aafZW9IsEy6pRbKU2ho2TZJBqu2JvAxoI5WJpBRDdbQm7Y0kHDopRvoavZ0VN6Gx6WyVaIXZp7Ho2NprD2aH2PRCb0fuesaeVjooukfh1oTpF0LwJXs7GnRfQ0Niwj7ENi2IRZs8KN+DFveF3BKNw/B72ITVE9lnQn6WC6Gui08LqjeYtyTonTobG6Wjq2TZcJ1iUeE5oo9vDzYMVKIomQRdHmGhqFK5hJ4ahODYhE3C6G5s72LCgdPZ6MYlcJbH9jcKXY16dMfeWeFGtjQfWxL6H3Bu6JB9nuh/Q4jwXQxiEqriPVGJemJqa6NwigzkKjhPRc7G6bKg1R9bEotGi+hvexsIN1wb0XzHZPcv7wtjx4WaH2ejRZoSHj/8QAJhEAAwADAAIDAAMBAQEBAQAAAAERECExIEEwUWFxobFQQJGBwf/aAAgBAgEBPxD+6/NeKXghCEsIQhYWEIQv+4xjwxjHl4fiyYfzazfFYQvjXwN/+S5Uh/ZfhcprwQsrSEhCwsIWELKQsIf/AFmPLYx4bw8seGPLGX/wP4Li/Nz4eiwvHhfhmEkP7L8l4rKGIQsLKwhZT8V/1nhjeWx4uKUuGyjw/gn/AJFlHcvwWaX4EI6c8vXxqQ/svC8ELCIJ+F0ITFhZQhCxRCE8J/8AXeHh4eH4NEINDy1hrzmVi/8Agub4c+G+VzS/N0XD+2xeVz3CynhMTE8XFKJlE8piFjpf+ox4Yx4Yx5Y8PDHl/DS/E3l4WL5rmL53yWEP4N5pcLGsLh/df+iJlYXh0TELFwmIWFhCELKELC/6qHhjHhjH4N5Y2N4bxc34l4XNL53zRflpWUuLC3z1leC4f3X/AL5rxQspYQsoWFhCwhCwhf8ATY8seGMeX4MbG8PDw83478q+K4vyTPvHM8+FcP7r8V8CYnhOYTExM6JiynhYomLwX/SY+YY8sY/C4YxjwyeT/wDTcL4ulPYsXHrLxTme5s8aXK4f23/vhfFeCELCwlnghPCEIQhCFhCf/SY+YYx4eWPxYxlGX/w1F/8AVpF+K4vhcXLxfRSibh/bf+57hYQvBYosJ4TELKwhCYnhMTF/1bkxjwx4Y8N4Y2PL+G/C8XZ7nz3N+SlmKW/BcUvrwWE9H99/75LCxfC5RcJiFhCwhMTE8JiYnnv/AEnvDGPDHliHh4eGPzfyQY0X/wAd+alL8NxfBcP7r/3PM88Fi5omUpSicEKJlExMTEJiZ+iExYX/AEGPLGPLWHhomINDQ8zD87hY553HvxvzX40POi+dL5Lh/df+5XhfC4pcfwLNyhCFhZQhaExCwmL/AJzHlsY8t4eH4MeWP4p4XyhCGjRplRTpT+f/AAr5H8FKfzhcP7r/AN8F8y8EIQsrCELCwv8ApPDGPweHh4eHB41lvNLm+F/8lKXxvxdOk8X4UvhBWKDKWisP7L/3Cwvgvin4IohMQsIQhCwhCFhC/wCax4Y8PDyxDzweXhjEQnhPCE+GYkPQ/C+SzPGjL4UpSHPgpSfZIVIv14Lh/df+5XhfBeSFhYQkJCWUhCQhYSELKF/zWPDwx4eGPDw8PxeF89+GC+SiH5XHClpfG4pTYksW8I2ReKkP7r/3MEvGE8teKEIXjcrKELC/5r8WPLeH5vyfwLNxs5m5ni/Fl+J+PfKizfo2TFI2SeLKbFw/uv8A3K+RFQmJ5ohMpcIuE8UWExMTLil/5Tw3ljGMY8PzeWLDxBj81l+N8oQeeY4MaMiNGkRPhc8F+Klxov0bGvKm2TwLh/df+/CvC5RcLKeEUTxcp4uUxCyv+S8N5pRsbHh4eHhZo2UpBseX8NxPlhBk6Qbiw0V/+DUcYx/hbb4UF+DRUVFysc8L6xvEWL4rh/df+5X/AIF4IQsLCysJ4QniiwmX/kPwbGx5Y8PDH4vEFhomJ8MzS5o8c8+3hqjoypP3CNuIZccId5ispSs2R/ZCImKUuNnRoiOeHvxeFw/uv/fl3mCwheCFhYWEIWE8ITE/BPC/4r8GMvmx+Dw8Mawv/JMT4O2zotY7wXsjsSiR9veIQixw7mEIQiIPDy/B+KOZS0f3X/v/AIL4LxQheSYsLCFhZX/Efi8PDwy5vi8PDwxed8r534bBdvFO4Yw9D7F9s7jh35b48yyeaekf33/vwJfCsLyQheKFhZQsXxX/AALi5pRspcNjZcUpSl8KUbLhuDZSlKXFKUt/8V+iD7aP4yxiU32EPLPCiITMyl48w0TmIQvnzKWj++/984czMd8EL4FjuU8UTxRPCZSlExYomX/10pSlxSlGxspRspRv6KUuLmlKN5eH/wCKfD3O7ZeIaoJv4z52tD38Dy8Ja6f22c8V40uacEy4pSlEy5JlKUomUTEyiZSlKJlEy4TKX/z0pSlKNlKNjeKXFLijZc3FKUuODw8b+OoqLSlEP4J4dsbEoTHESIHiUhGdJ8vS8di+j+Tng8KQ/vv/AHxnjc6LilKUuFKUpSlKUQpSlExPBMpSlKUpRMpSlL/4aUZc0pSlG8tlw3l/M0Twg8zygo6SobQTdY1fBtLptwr+iF0Tq1hLEou6TE8An/0xMQhPCYhCE8e1iYhPgguH9l/6MgvBD8b57yi4XknhZohMTxS4TKJ4pS4pcr4OFxcUuaUuGxsuX4MeHl68X5shBZa8IQmUmx+gjb3mGyMm6NNaDiVCT6+idITG3xCW4QVGnz45oQnjCEIQh2iEJ5pPhC+st0KbaovpP7r/ANyjvnPPvxoWELKwsp4onmiZcUuaXFzSlxcUvhRsuaN4eXh4Y/GYg0QmIQhCYZCDRCEGsIQhCENj6JPBkEFf0OYTf0QbPbGol+irh0j6Ij8hhotDtzKkNr0VGno4QS8OqiGHN6DURv0R/RfUFyPq2M42MvguYmNCbxDO2ewxcSEiwv3P91/6QnlCE8ITyhBLEz3CwhZWFlCwsLCeE/C+FKUpS/HMNDi6fofsP6ROTfcJ/YegHPh+Y/oQlPext4hyUSkCMKXlX8cX8Cfon6F71gt7E3jK2iEIQhCEJmEILwNVov6KJeiTN+xvXK/cKkjXvCVNfZJzw4nTMH4D20z8MfqE3tk/YhINEJo/gleEiI4zTGx1o/ERpe0hJL0LeU9nSndiKf3X/uFmeUJ5QmIJEzCEJhKkxCeCwl5LyXyUh7Gv0Gv0Gr0H9AaQ0rp9sHEDcG32G223iEJ4P4qX4bhfYL3BN7QndRb2J3sTOPEGsJPpDZwo+i2jR8UTKcxRyf5xcUqBCZKi3inBi1Z4WEIYjg0TNGLpVzHBCwoXD8H0uKJwXBv/AKv/AE7iEJ4zExCEITM+Giwn4LCeEy+FKUpSlzR9zGAjxj9CY/qH6Ehv4xv6G3rDZ1m/ZMTEJmeHfnfg/JeVxT2S9iTxj7mIWKOO4iidxSlH/rFKUasLhdlxfOSwnhRncSH8HRQfcVkXo2J/AjZT+cJign/1f+5mZ4zExCZnwTMEheNRC02NHWQ6xN4z9hfcfofoKsp+guCYlfsg6YS4bG8AH0MNEIJEIQhCEIQnlPOfDfL887ljz0c8dFKXEbcTKJlKUR//AGXFODFcLsuxb0b0LTXAWF0dHTvhacNLZ0jYnDrGzgh/guFKLHBDeWfmKLh/Zf8AovlhCE9FJVouI/op6J9D8CJ6GGF+h/oj7SPlGiThH9j0OnRseHhYWfRSkubieCKVlKyQVFXwzFvwIeZh/IspfE8aoPuJlKJiE4Ol/uJzBBO5FOpTYhuscPQOJcJlpYWluNvFhS/RdFQmXDRwTHFj9HjomWdEx7OYTHsJ+z+E/RD/ACPWfwYv4D9BP9i+7J+xI68/EX0i5ET7GmDWHhj8HiM4P8IPmGOo2yUmb4ouaUpRPLZTvhcXDKUVlYwQVPC87leU+TngvDRM8DuUomVFjKJ0bf8AkpRNCOBUymjwZ0NGbJsdyaoWnoTKLZTh7FWczZ4U6aWP00xjvoSf1n2PhwBgW9DZCc7DdKhspfsbKNwrxS7Kij2UtRJiYaxCERo0aLjYyDHjK4Gj0Q6NSe0JsGqRDQNYNeCKLCKJnfFiKb+JlKRXvGCCovlvxhBL4XzyXg3jgdi+CZsJnQsLvHsbqkLTqVwT2hthPTxtYaP5FrHrNE36wTNjTR3ImKibpoJOIoYImhuITY0moUWQ2pBPI19BI9CSIjsN4KbOArqI2X7GngxH2JIiIQeNQ4UpS5exjRCeO2NGiSTQ0k6PeINJkQkGqRaNjG8XD8Li4paUuKXy55PxeVilZSlKUqZSn7jXxLnws4HTx0UTG2KLFPT+S0SGZcQjexWEyRwpvBLYl9CxPUxEn8hC6ElG0SXYU1BsfBJwaY0Xo1CNCQlOnThfwTFpoehUSY2yJLEJoROsNU2JSEBKC+4xPRVG5opWUrwtw1hsuG2bxRtlY6OlZsVbHDTYqSCRBsb1oaLBvDZB/eGP5Lil8L8XPhh6+FkzMIQ6xZssoobEZsaYx4uhI1Q6DVEUNuQpiY9DQLTIjfBzcE1E1g3QJvZV7EqpErbEgMKJ4W1CopC4KdZI6QScNkI+j2hfybCCRqRHNCWCX0Rt3EojphoSQj9NshVEl7IdwgPNKJjg1RY6UpSjeKXWGUY3h4ZopcJOjTQ40axi0hLhSjY0ZcvLOjzPG4fwI4XFLmlxZ8dxRJGhjOGyC1lU0Jlomd0RiEt6Gj7GxHseIRSPKK2DRqFhINvRKPuh82JJqCU5jbYmJstWF9DdUEINDODGh0osIgkNJYlFWjZW2JDRNi/Rl6OnDR9jFXsijCXSQ0pD1g0dxhEtTHb8F8GJDcRtCsTGz+MbxaUbKPYpS1j5h2xFmqSaxKhwRDRB6H+DZCvomNjIUo/Dub4XwuVi5ubjeH5aKJ0b9YuzvhcSkwvBBIggghfovtD/AAT2UlINQ2Rpo2Z9kNum2yNbFfYjEfTbUPoxNCQoKkqhqWCbE/sTgmK2cDEt7ODQpMJibhsm9j6BwJHpEvpF0M3bFRUP+gUbMY2N1tkfYrWj+8XuYmRTf2Nm2Kuirgnga+jUEH5PB5ZLaLBjKXFLBiNjcG9jZRMbR6AzWxjehfobKX0bGMox7Ib4NxjKhjH5tn8FpcLDwiiExsRdfBRu5oiNfaHoR+5mUhZgni4SIP8ADaWy6FSi6xTEmsS7NhIhacOiuC/RNXhD4JCCUIOkNSISoklsUeEhA/oWfQixia6GaVQn7Y3aLFaIdxmm0LanuBiKKxIuCEhMnREjEerG2CaehhDfQpWD3G7xSoSbQkkdKWMTZSzeD28zEHmnobZ1BiZ6otY4VM0Uk3i+Gxu6wth1hLbRcPDGx/Yy4bw3Bulaw3CjdzTZcdLPBDEUWi44PCY2ey535JuBt5T+youLhXwTxSYSF+G0baILWEWcF9sW8Fo5j8IbIfgihoiIb0SkP4E0i7w/waa4P2IppYku2P6H2ikLbbIKJ1rhqDUDTguwuxVoaj4OtaQ/2INiQbp9jQrbBUTb6LQkOUqRCdF7CEhGxIaEmUbI/RfzybGMvobyxtA204MSmyCZqsb9Q0MkHYSkNpsYvoTYiG0WDKMbHoX2P7xcM500yMaHjjw0s0b8+k8N5azcXxmGy49E+z8GcKQg9CysT6PRKQenoW+iQhK6J6LNHrZ60JtI2Y0hucFTJSUJ6hZs77LvDQlCojhPMKDexp8GmlsSBMuDTSoiht7LbeD8hL7JS0zQECSSG3gbSEfoWkYoeW4J0TXD2RDfpE9CcpCbWiNnR0KFi7Ejo0IdEiEy9nB4g9DzRs5E1GJQ/BCTWC+CNFw6tDwIY9ixHSHvLWPzLyy3DHofg1hv4aUp3Ceb4L6JMvD2PCELD6NC2cLoRsV6OorxfWFCP0/ge9iVFtQhCG/rEom1piYg2Pgo4KjwP6F01RRGmLpKJfsSCWzgmWEDa9i0PYlRONCo0N3QnDRskJs4PaIUMaTYoMNoegmyH4VlEFs6o1NolEiGPDGiE4WIa4hCj0VnvyYzpPZbj0NISILHC4tGcqQ1uGw1CzR7WSPHM9Ho/gYnRsdGbEiEGkTEGPwX6Ue/GeEhPBlzwYmU7jTQyliwmht+hrCIISEOEolsgkQ9CNBVlFMag+CnBKDWiEhESiIJJlLmDfokvYoNP0I2Jeh0RoeiUhsJBITPFJ8KxYDV2sEwkFOieEMTQtiZsYL7YneiRb6JBIxIacKQkg6Ko2nsTo6DhUL2YIlJok5jWxX3jprF8NkGqQbmHDw1hO4ex6FRI5waaYleDhomFcsdG/Z7Eq0IYlGPY2SZcGIP6L6J4vRceyC6PHfBbzrD8FwYxFPZwuPRBoiSEyehJlEdENlINC0dJ6HpoS0JEdJ6EJhIQ02MgyUjswjmBUXRr6EQV4xLZ0W+HcGjx5o2IFKehCDZMWxBDNJshcGm1RpoQm7BUEyp9G2IJGUt4K8E9bE6cHEJ0uy0dG2hN+zpVF6DYzU9sTIWmM/RTK+x6e8Ri5ljQezgx/RwZpsYxaEK2e6Qobmxsti+iRBobTHiD/B8PwdQ0N/RzDHopR88IPWEOFyhs74+/BoVHMUUFo6MbQmUXRHXnqJSDKQjEy+sdIL7EGJTQSiwglRqCJsS+xcGmEJoS2NCVIc4NEdGuDU4TCUFlEo0Y2mismxUXRODLHoc8HqNJOEoa9EGkao2/Qp0J7cOxsWhLRxG26Jij6RdNMk4T2NbHt0ZtaFPRalCVGq4xc0RaL8JdEZqnRnrLG8Pez+RrdHtUNf0Jv2KW4jpo2OJaNhIRNRlHRqOFnRD2N4Z/OE9m3DTZobZr0NGjQ96Y0NXR7g0ijHiHCIein8kzPZ+nR6zc8H9n8+FOkRNCGJEQkhkEiDWhIuyXBorohht+ht0ilF+hoRfvCo/QhFGKNlok6JEgtiU2NQSL9ENkdC2h6Ea6VUUOCZSU4g4ehIgzaLEKsgxJ8KLp1R9HWzh1iEyUqewv0gVFrG4N6G9DpwLRfvEIINUS9k9l+hp8CQiEvZMP6LBMrQ2hiBabZRujfohpwa9CN7F2eiKujGxcEj3hE2JGJJZmhqHSD0MarHoQg9YSSHSbpcfg/RjWGfpBzGjoywp3C4PHCePTZRkuEiMQ1RIhCYQ/oSGiJGhLHGUTPZL0itGk0IXDcaT2UDRwb2NG+yH2QSdNhIaPQgho54exwgYuFZ0TJsg1Fs4Lg1WWDcGJhKsa2P3RBbZWhwMKt4NUTWiCHuJ2Q6J+hncQXSRbEqImxo6xJJjRNC10arvhvDTEHUQ2YyEIPpaegTehphKGwxCQTfscF9i0U9nR6VGetC0x4pQxo7hnRsZB4bSLcN5bHhotyhJEGTE8YI6LmITDIIkOkjwxBibxKT9NodK0Ig07RoV6QnSPQ1C2hP08EkaSw0qPfBtMcQ6fBQW8N9FexQVMbUguEEhIgvodEJBaEP6DG4aIJsQgwn0aaEjFPCQaGnTYs1zqRhiaIdGuxehttiLBb2KEglXSEHsJEIQ7zMIyl8afo2UtN0E2bGpBHs4S9Gh3Boh3SIy0UEMg9LQtoaQmPDUEtbH0mstDPsNlmyoesJPHsiW8PhJj9OiWiQhCEITMxBQnhB4jEoJDITDwSYomUQTHLwhvh9RLJ+xL9lrgb3UxFPQNzUs2DX6JLaGVVxG+Nkw0zYmQmPaItwdXhLmxpEIQibI1iYcK8TCVIIEJoSESYNE2SG5NEQww0SNQS0aI/A3oTKIkhBqn75wQyUmHh42aGiaIPRYbCDSJ6OISvT2YIT7GPRGyQUdGkP6NlG7o9jRCH8mkaJ7GvY02NMdGx7GiIa+sJsnoZ0axDTINwSqEPKzcfuPY0TwWjXcUlFiDWYPY2tQmuzrZA8N9RYlBKbxpkRDEpwjJhul1s0yiLH0CRuEPQ2utDW1iEGOCaZJT7ULPmicS2K+CFCo0NDhSHCaIJMjEhbEjpPQt6O8H3MxKQ6NQSND10QsE0tC1gmI6L9yiE1fHmJhsgbOFxujRwX2W4NC5BoSGlwo9miexjRIQn2OEP0JNEIbThoZEPRD+SpiR0Y1rB7GQag0xQNDRzQyERCNDVEiFEe8TEZISH7iCTmILWIQ2EhCxPZEPpPQ9dHoS9nWb9FgmhKi0RMSgxBo2hRHBKGmTBaIyEjwmd4QSDobLEPSSNdCqvgmibDRsa0xqcErTY+tMSMaMRF0Vkb2KvuIJClw1OEokPhMrCSJh7wdDstqit0RDnRCcE7hZnjcUf0LsbH9CrpaX6NHg64LSGmxJp4eZ6Fh/Q9HR/RNCE9FHD2Q24UkWkdG9jZxFLRv2P7NBqjElB/WGvoS9D1hdjG4LYkPOzq8ODs0cFGXZ3hSrCwgk+kaw2JEhBI9E+sVFtwctDZMX7FeiXp/JoJ0c44I0tmiIaTw0OipBDREzngjhzZ0nvCg1exutoixGhTg6aZvtHSNJODmUa6bNFsfRJCIS2JC2cR/GNidEOzQqLH6fpUfxh7RsWyB76KTGnqCqRfsbRCiLsvjRYlwi2JaNDYa+xtjrJR6ItjuG9D4dh6wzRMNaIPZUtMUfMTBDdITZBjgg0mozQa+h6EhtLo2uja9DRH6PooPolQn6ZsMgkHpCX2IhRcLHUUZIWuYtGGoJCVIQn3iEEiCxCbGMa9FNj9DEq4UWiaJ6WCxwiHrhBbEtHRGx4RCQn2M4UTOoglhpPolXMUWipK+iGmi8mqhPQvZ7AapI6xa0JQ9C2QSuEM/gQ1hLdHUX7PRKLYyGkxIhNjrBh6QlHmiapS4WFlEDXT0SvYlBtM0Fvgj3CbFootoTSNCah0Zw1jQmh1saolENj5o9kFsg1D+R7OkhBkE6iZRnfZjUZQRzMtxCpbHynWP9NcEhDrxNCEJoTKQ1l/JNjSXDQ1CiEQmyQlw/gRBLWYiaLYvqNMkwyVUSmyVCOoRazQ9H6L6YkJRiGfotcLhpIX4PeP5LhQlJhpQaXBhHutMRTY922hq1ogJiehHdCeOHRfQzpPYsPYxiGxext4lIJUhNCQ1SJoQbIWu44e/BCfhEfyexPZSoaInw4P7Ju51BG+iY+DZ/I2hI20JRL7HoepBzpnuklg0PWxOoYkdEozfBWiGtdipI9Gi0MINboWmhejZSdh9paceF+kohqnBdIT2dI+hNPhIQdeyCEuyUQZ6Gn6IQcY1SRiFiD4UmLvOhL2a9F3CCSQ8CR7g9D+iNaEmtDHoUZFSC2QWNDEM4Q6SI/crC0TMGjUNAQh7Y9wEe4gml0aWYKidFruWrtCV2JEFhDYlj9ELuIIWiELvMxDaNM4Rti0XxWPePxjQ4TWjR4JoXD9INQRxjF+j1tC2Jpwa0DZY6qUr8Ga0cFU2fyd2MrCEZNjQpOmhDdhLVQ/QJ9BQtjQvqUdSFdNdo4M+glQkxGKjTYlINRaNkpBSg/gNwaogkRCGdDWDRIT6EhCFSEH9+C3somvWGR+jhvp0qG6NV02RR/o3sp3bElCEgqxIImEyHsez8EL6OHWd2N4X1mYuJRaZNMbbuip6Eq2hf5hiV9i+nin9C30kFGNODfZBF2eso/ggodN8ws9ZPGCQxBKHDgrm43juYQhPsSgl0kINYY/sTUEqhJos0xwTiEGi0XtwkTovsSE+hpN7J6F9EP0dp6QmeyaEk9jRNj4Ij8JvZRQpaErrKPTEoNqDL2wkGyTYsbwOihanRKkzgSOEhKIZCCWDwRvaFWhoyjexvH8j+xhtM2tIVS2J0f0EzoajoR/BIOjvsmxK9ElwkOY4JeyHvEWGn7EmhK7Ix4SFofwJkJoSHYImJoSsfB+oSV/0aIELQ20Jr0JRTtiSNEfZHonoaYTDV2NJkIJCwkTZ6NCaQsdFHzx4QhMQmeiWEUMg20PMw1o0xr2NexqjUJFspoh+k06P5Hos0N1tFpCbHvQhGNREHvgqWiNcGrwsa9MSqCSSINTZGtlHo9jRDXsUlBp3Q19lJtCX3ieyDRNYg2NsmyBacEjjNiHaSkEsiekIjmiERp7E46zbZbo4XBXEKlKd4QbjE3ogURW9E2cHvH6sGp0WsGUS9kISCTp/Bwbon6NUc4a9CHRKEyhYR0/Bx40On6DjSEUF7IIKW2zljTrEJUamxbRMTQS9DZcGvUODQsWno4SCRaFhC+yXHceiXEvjCEJ4so/oVFh6y0Phfs4QT0M1Tg/0ckEppEI3oWiW02CezvDmyaNwaoyC6CEhn2HYoEmsN6GOI/T0JL2e9iThV0olRyiVQ0QlGho3Jei+hV0S0JMVENCQkRHqjNiEK+httjOiRvZEhouGyEtGzhGJNsWhp+h/RtzFSDUY0z+Rxw2JUShCE9CEhvGh/BDY1s3cTZPZKSvZMJ3Q1o2xYcpPRCCWhETIuEMyutiiUZGjRotIi7rYhRfY/Y1NRjiRsZrg3UMTYh/ZpCGayj343WEaxD0eiYZCYeIhj08fhunMbKEEGSk2QY19kINC0RZJnSREGrpDGtREcYlEhc2VPglBnrE0KweiaNGNDSkRsJXBoV6HHRaUF+CWofQUH6J+E3BhCRiaXRfY/o2JE9YieG3Rs0l+j3BbYjEuqV0Qrehv0sMSJoVMaSXBWqLTp+spXLiNi+mSk3BfQQWJhfbNtk+hfR6lGQapoaSZRU4UUH84UxKbGSkwl9jWxpPon0OIljbGsSYtliy4Pl+yCw0o0AolRME5xjRIRWwqEspqYfDgmTKOeNxKIb8N5gxx6xzZD8Nj8HhkGiIg0mexBoaEieyQl0RvhBq7Iz7CX2T6EezGdOdINQar3htDJRpomtD9sSH0Y/Q0UGT4Qg0hrH8CJCXEqSEyC0L6ITCG+LsK+xQNmb9Cat9wSjKbpTehOlYvqNoWa9jY2LfBLVJCQW+HR1CN9N8wvoSJUKkLkLMRYnCbIpR72yLiUhIQ17EsJfRw2INCWjhCHRHoMdQ9Y1NNC4Tii0hRT2Qm1sdRBM0xo0JrUJWJESbbFRbJFsgtssK4NtOC2aEn4IWL4ejng/HrokNCG8cPWLsm/B6Eexn6NEpCIgomiQmNDrLw1FTvRiE2NbGibJuDR+H4cNhqOFXSNsT2RwkO6Id0PQkHtCsqVCUqLqix+4lNiUmKkOCbYSnBOODqJNQyYyehSNE6LlHCG6NRv6OjlErsqwcLRvVEm+iojRadYSLR6FwS3DRid6PSF9Cqk9kE5omj1hmwts0JiVEOqkgtK4usJGxbHpm5TaJSHdB0NMb6PX4PwYxsXyexWaY3Hs/IiyCpKiUE4J7HW9kYwvwWkNEhN+H54LCxRoXD0IWxsWP/xAAqEAEAAgICAgICAQUBAQEBAAABABEhMUFRYXEQgZGhsSDB0eHw8VBAMP/aAAgBAQABPxA3/wB+UMHwHUGYQM3BAqXMECfRCAxBcECoGJjAuYEEIMw18ENw+dP/AK7r+jSbI/FAZpHU5i2fDt+FjGNRgq4/Bam2ZREXqOYuJZLjv5cnw6l/DC1Fiy6ixGL8DLly8Yi1G2XL3LtqLE18dzc+vl3qLccxPuJc3EuafCRojn4ZXxUQnmJWYsYuZb6CGv8Aly+AYxD5KyAZ4oZQmMQHUFwCCBKIMXDMCCBUr6QxBB8B8BT/APbdf0Mfh1GO4qjgjqLRFbK+DT4GPyByixYxcuKLE2nqKxjLxLJFai4IjWZmpfxx1Lj8/cuXHMzoixnucR3qaSr2zTMfc18aj8Vz8MSyV9RJVx5+FLjfwk4lZ1Elx+DBetxGU2GiH/t5YYGCekFwMTOekrU0l9QJvA8w1F8AxDcGvglN/FGH9A//AG1z83Xwvw4Rai0RzuLUojaMYqis38JmnwYwWQYInwxxj4RmZmN/CXKfr4Uxj8PiwykfyjFBuVNzmXRU0SpVt8RzK+46ZWLlX9RDxP18MW454iJFiSsRialbjpzMRPjiMdx38LHUX4Kb1Mk+pkf/AG8o4NERi4+XxDTiLUUMR/CiislxRWQiuE0il/Aafgag3D+gf/supl6jr4cwROYLJsqJEsqDMS4kSBJVPwwTJHCMOUwxlyjCRMR9xPESJ8J8OYseYxxxFOIsZ6i8Ri1uNVGXLr4XGcy4tQeeJssW5cuXVxYsU4l5i5ZfMuLmN7lxcy+ZuX4l58RemXFqJzF7lsyjZKcGiOl2/wB9F8B7llMQ1AWYVFF8GSDU0TVLPgIGyDUybhAkKQgpMMG5dQbgw+R/+s7+XM18hHXwsWMEdx9RmEdznfwzaMYxYvEYW46ikaixYx1DTLixf1EYlofhcWXNTccHwrFvUyxOdfF5qMPhfEQ53KF3uJi/h1PMcxq44vuLHJHxufc5eoxm4xzmOok1qV3KuJEqJceYq9BHXV/fRfApSU3FD5APwYJtHcXmXFncSQz8C/Ag6+DAr18BzNw+dv8A6zv5dTUv4ymkWO5cWZvE6YsCpkiy4wm/gbRhlWYq/hajLCrFYuIsv4silNxYh4iLjwik6Rcy4r8jaW/D4+blRIniV3AjuApHFRiqlSszaUSkPETqfme4h3EGVcSJXw8yoxqM3uNGJF+AgXF/7okQlkt3KvgLQCBiAngxAlIIPgPgQIbhhhkmvxhA+Dfxz8kv/wCo6+X4WvhYsxloxvmOpdxjFubYnwbGJHMSJiYQY3ma3GLGMWPUrEZuLHMTqPccSoxlMSJ8eamplEplSq+X45m/i52RuW2Jb1qOZti5qO9Rz5l5+Nu/hlefimajqOfj0i76ixYttO4zpcEv/wB+0UEwPMGI50g+oYmUBFUEr4BIEG4HMRCxuDn4BuLuGINxfJdMG4Mv5HP/ANc7+NvhRHw4cRYx+YmYykdy8/BnhH8R3UYIkTCwSriQRImImJqO5VRqLH8Rb1OZd/0LNx+VlfcRqcRJxHPHyzZOO4uJecznUpyjuOopqXqWRcdxzr4vvMWfc+443FuMY7it9TRNEcRX8B0aOZ/1e0pcdRBBRPcSwYMf5ggVgv4EMwYbhxBnxAIfEhXwGoofA/A2/JiDf/1jz/QGYES5e45+b5+THD8OJhGMWKosYtxRcxYvcWmXF+FzF/MXMXPxcuo5jGOpfUZsmSe49/CsTW5uG41qXLiyriXKCEfxKlXEzWIixIipTPUrxHwiRPio4mDrMVHwlYziU/UTZKiZ1P0CL/l5QErAhASlQqFRg3BN/AoMGKK/mMGDUZLuDKXBg8xTcMQbIN/0Dn/6bv57+HfwppHUvP8AQH5L8O2MvHDHXwGJEZUS7iWRLguJGJUY5uXGI3fEStczUqZ0ESiVEuVUfKVKbiuJbmNJdyy2O0vLx8oQ4SsTCV38EfcYZyJVGJUQZZqOPmftEwxO8SsRJWZVsTn4TERqIxyiZxEcsBo4IuP/ANUddXCkMofSLz8BlAVMFSniWcw+IcJRD4FwghRVBuXFBzBg9QgbhiDcGX8jX/0X+h1NR+MMfDScfC45jv40iw/EZWIG4xGMTEETEoJUqIngjD4xlIxl8FQsR8fiw4RJUrPyqVzEtlXKjExKlRJWNRIncaeJdxlTEZuJE3HLGxjHZ3KxmVlvUqOIzzHe4vcUI838O74l58RU5n65H/28osfIInESwXuJBg1MhnEPkAyiEkmUK/CR0M7YZwdTyTZBig3NZhn1Bv8AoNf/AEzEjqa+GEiRp6iXEqOMSVEuCInNRggI11KLiE1GozEZi48xYootsWiNy5c7i3HB5jF8Rj+/h+OfjcqVK+EiaiSqJU7bjqo4pm5fw38N/czUqWlc8xyj+Y2NT1+4/lGkrcTMSJ8EqJTNM8S3TLswfmb/AKHEf/Xyl3FQamT4F8BHS4NxWbg1CP8A1haUkFC0MIfAHGIoMHEUUGoNwcQceYvga9Qah8jUM/8Az1x/QvEcE23/AEBjlfm2Y7jiLFuWnHn4S50RImYkXHwiuoqKloqoriPnGWfaDGkRKlRBcxCIXEES3iNMa/ME+GvgTqL8XLxFzL/MVI+hGXTqOWO4zmLuVRuKa/cruO5USvUcseIxmo+5xKzOZj4sSAcs6d9J+JXJl1o/EwAUHiE0miKv+PKZpyhFBfMHEGG4fAUIPziRLxEgsFZpDMJlA1uWgQfATlDcIanPwa/oH/5y5jv55jEh8MfgB8NRLgpjUdRqopGa38Kpki37ixdy45TBLlxZctJcVcuNxWZjmZ18Ln+0TMC5iMRlMzKlSmVO4nwnyJe4r7nOVTHhAZTfwfCMZRw18FfF5RvMY4RTHWPnr4eUdr6MmVxe7LE7D7BidSjwLxLDGen9TW2iXX/HlAJTC2oMWe5aoLYFQAgQqFQoiIiCRHcBCBg3FT8gMUNTiWhiHEI6isir+g3/APPd/wBG4tE4l4juKtfK8fDqL5EYx+MoriIxIkq9Rl8I/A0Y+EfgNJWOWJtBHL4VUYpGPGM46I3YzcjSOHwYp8KlTtE8QLiIiUMSo2Y+JtxE9SrGOZX1ElYjDqbxKpghFoDuK2R24I7LXoIBQDxDbAeYrZ83BHg7/nM0RffMS8z9An/H7QY8xYg4g/XwKWxMCHwH4DcCpvmCekDEECoFwUVAYL6iQMwPgC8SoKIwUQL/AKT/AOc/Lr5bjHNxjqMfh1EiU/J+B+/iswjHn4qJcYxqVOiMfESJcwmmMQiVKJuVmNHuPxuVMDK+KsZWJVRcxxL/ADLrUdSsbjiVzKiy7jLjie41N/DmNTiLeZbFRaN0S1Vuj/KJuA8ZYtYV3lDbQPMUs/k4I6oev84Pure3LHE/v8M/QJf/AMeUvlUaDixbIP4DyxBhAsBCcRGoBxKQHXwPXwIY+F8D4DcMMuCxis/qH/5q1/Q6Phys1FHTFixBFo+FojH4wupbn4DUWMVm01H4YkYxYxiTHqMq8ymVUc5iQ3E8TnJHPyu/hcdRubI+rjOYtwa+afjiLGOJvzOJ+/jXMIi7gRxH6E0rPoXL4A85ZV3X5Y/EUqz0LnOA7dR6d0a/cTsM9uWNKn4RIKiBaA8xuw9JGrQ+csXJqOCHj/8AdNIp4Q1MIJeW5hiBAhiBXPwpUGDcGDBh4lkIMHqWQYNwYu4MGEFGDZCH9A//AC1i3/Q6+NoR3GPwW4/D5juO/hZQi/iGmPw0wZjuOfhm4gx8fCwTcc1EjESOInESVcTESVEr5r8yogLWjuNe7N/dP6ikMSCVAbKPEGLfwH7fxzFXx3Or9n4Wtro2w/F1/iFbsI3JEVpmqwbgph5gfapPxKiMS9zcriMWlfmVUSVKmdQPcbfxGJW4HgtgPP6W/wBS9B9wolbfRLZZt7WPxBaAHj4fMdQAtQPMW0WvC5/KSjhoHQqDryd5Q1GW+onFf/dE1O0HwIoq1qDZDEGXTFmaIOYQoL8Ch8Aa+AaPguWQYN5iig3FBshuoQmn+gT/AOUf6L/EW/jf4d/DqKLcdxii+GkUWLj5YWLFjj4tcfDcTM1MxGJZKZaJEZfMUy8aRjT+l+iA4z47+F59jpcTJzvU8VQB/BKbK0bUYDOLTg7IFfKNoLEepWlbFXcL9B+4wa3LC+uefLRzE9Qz+UZ2v4KIiKUKEWRq9blBVESJNRlT+IzZA9sQwC/VRJVH7f1K/tmECyK7csvcnoVPI9lwHA9ES5tHG+JhEX4Zm/pK/mPF7DcX2V4BKM5PnMoFVUbYm05OJT4P0iU63++lYMLr1E1BiWhu7xDj4O4IbgqG/kMfAh+5X4OodQz8YPyDTFDcGmDXxp8DZ/Qb/wDkFqLf9G4t/C1FuXmO5mJBHcSOonySJEgi2fFROoxQRJ6iSpWYhHONTUYTETPiB8J9xmtMSo5lZmpgIlfDqB3AKo245/7mVErZKqMBc0yw5/BgCJTikmpakZDd4XPRxyQbIgEjVJtjReUwQSBxCsP4vJ5szxD7ghiAMUC65oiHlQTofX+4kor+mZ6T0M4gfj/cp6f3Qdta6CKOw4f8IBr84awfUaOYDYPbEeP1HzPpRV4brFToJ7Zb/YXFtp6xFbp9lwOoV4iF+ImYJUt1BGO6iVE3P1p/x/L4g6mGauZQL+AIEsINwKgLA4xBieDECBCEK+fSDA1BgVFCFXBF+CoYJdkGsfA0y7/oGpf/AMZb/pX4WorU6+GBcET4E/MqolQWxK+EI4iR+H4eYLYypVTia+GVcTFRVxMziVZKjFiZSs4jSbSpU5RJouQD0ZKmd1HcCKCIGPHTliiT5Wj/ANuOhHLttowPCdinmEgbwWugd6DgztglpXpidhDq2VR4v4lfE+pQ44imwibsfiPTPUX4/cet/MbtfuUuk/8AOgXD8T0lYiEYSJzElZlNxIn/ABPSMJRBFbIj9xEh/FP+r5Q3B8CZcQ9WzUUH4XTMMUIL3E6hCiEIYg3DEyg4r4cRPcG4bhuENy8QckGKEGpX9J/8dcdxwf0K64i17+FhHMW45j8LjU5jGqjOYsSvi4pLMx1uXMVv5u4/A4RhfEuLLhiIly4sWpi4pcvEAWyjaxu2dNwwQRaxHbHSFBjEWIbXWMpuE8YpT+0rbcvbGXUWXZUusfuLF/EXHUu5zLuXWpcuLUUlhLi5np8MX8LBii3qXuNuYumIn6RKv+nKYIIQQAguCBA6hD4D8DDcOJpxLQa+Am5p1AhuDBcIbhOYQcQxCaQ+BuLX9A//AAmLf9Nxb+MPcbePheYsa8xlv8HKKj8F+DDLfUWWSnwN7j8V0Rw+NYw5R8/i7ZmMcpSR+N/P5FMVUWXmbTJWTKavfBeIu812CcGLinGT3KMrb3GHW4Zjb0S2XsYA087wyjqApOT0kGLHG8zLdZg7ixl0fDdR+buXLuLcWL+GMUDUA4O/zFxfHwjH9R1G68ymKlY3EQxKzifkjQg+oQ/9PKYcS0IJYQMzB8K1DM2YlEMrhmCC/gxAgQ3DUII+JtMGDjMVRQagwbgwgagy4N/ApBvfxfzdQYN//tYW/wCjmKEW/hpGFixYwywwwtTGN4qxajCxxOX4WLFzHJ8alm4sxdRY0l37+Fp+DtFl8y8VGJ/QTfwgZlbf7kAMR6LeiMm+QjvJADx8BtHgw75gRiOFyv2P7znWzLjUS4zWYlsXEb+XUT8RJipVMfhLYx3qAnZRLxiVqM+puama+KlPUTmOEco0jc2uoM9f+rAEArUAxAgqq4gkNQYMEIdICAYCHhDCFpcJJIJIGvMJIJMoLuEkGE+2F4RlBgwpCLlpLnr+pT/9Jb/ocfF9S7+HjLRixbi3GGG0WLH4tu4vwXUtFqKl38hCJFlVGcx3G7j5jfcSaioq4Iwy4cQpQhuxIa3rLFhOCFagfmkoqmupsWMDlXRqPRDTiEHpeGJX3EvxEhlMoxTZnRg7YVzt7Yoq29Q8RKQVKqkcrun+0aVM6FP3APPliTWIk5MLdXt/BTKj4RziQwllqbfDyhlGar4Ph8G85YiD4oV/j+n82bRymPx01GXnGk67UVf8OUIwQbhT4TGEknliAqEFYCA7hJ5w+DSVuGEIDDXMIMoSSY7gYecJBAwrBy2EkHwEGEHzL7lkv+kYMv8A/Dctm/6LhcUCXfxcW2ota+NkX4Y/Kxjv4S4+NfLH1DEyiUEcxFyhxET5S2MJE+onwTiPVYkShVtfdykYzyy/S+ZYQDGGIU8ALV0HcCzUC2B499sFhVmInDScTWyvMMmKZUZXVtX6g2XWKpNmag7eBe9PzMmPU2VlyWSzJ3DiWdv4gTRFDaRLjI8xyGsBAC+OIDhMIS/ALX/VP8wPGl+qf2mEYRlRpG0bR4Ssy+HP4sfnN/Exl4RS1Wzn1KmliYSbRrNPi1PcalRvPGPw8qI4yrAMdxQV/wDVB1uL7gr3uWOWDxBXBfcHEWC1D2g1CLqCwaiwgbINQYeUGXXqClwYrJdRRQeYrhSHSDBgwYNQYP5g9wal/fxdQz/WMM//ANLqLLx/Vv4XPzeYsxcfCyyJH4dxjj4McP8AQxg/OuZv4eY5+CNxIkYlRsRipgysQQgKyXTv2QRdyiQtNpdBp3xHscAvSFh7eWVhQe0bZy8zYCPuAsV9xTaHqI2cCZzVxKYoAWS4eT9kVUmW/BXu4AwKsvQP7+ZgUMDHgnm/BNs2woKUh1GvYwRQOKu5o9BYAxTn2lOmbI1PW42nLU7nozueOPAxNdzLzGwcE/vS+9H8AmcYvN5cjDn8bTxgV+if5RS8KRgesf0NIWyszlblOwMDxBEUAoOI5xXwv1GFzHiJhHtKCZyasKUXotjJQxieV4PZcbO03gzusHUGFtNGTymX8x45Sti17l3/AH5QgQyxCKqBAzB4YdNSiDxT8BiGfmmGpxC8wzBOJcPgQ38EIamnwqiuDmXUGDBmcS7g1ueYr9f0K/qGDL+Fpg38rQYsti3/AE6m/hai38s0fFYjGe4kYnyYxIkp+EzEjaYS/ESWJSS3qJK+D+MXcYXUtKiXH5bchlVqTkmHpUmft84CV9Rhs6dMwGcV3BegHJxDRqAFa4oZZxvKx9qRYaIP5So9bCDK1ivF2oXiPDhRUfu2K7yhTHIBFsZKwI+7RQxu9tzQMQD4EJtRrMBuXAGXzNsCeJTSjncWWKDNjqGyWwcj7mAXFs2KcWu4Yj6gA3neH9xT0lkBTt5SGIzgxcVQ9kpX8XdDItVQ8x21hbQ33HkXRhw3h6+L8VOpWV/MZllN0Di7ZjeUs1d6IijAqqVbvGSIllCyNtqSvFx40B1IpcZnnhxh8Mv85R/JIIADEHP4XTdRQhXkXyi7GZN7vY+pXipILTnYzwwtkU7DsjRzHGJRIyqghwKKo9b5glYK/wCU0H7h/q4Kv0W/uUVEGIHyOu4SG21i62qYVXzZTuggORruJTn7lur/AET/AJXlEhNMPGWhJBjUKkPgIohA2GcOFXKhBJAVAgQQgQKhAxAqBMPjyhjUGpcGD4g0wann4GpTNvPxUGviv67Zdwalv/8AJmJ5lI7g7A9z/wBSJf40RaRekwl1ha68vRBm8PUb4Dp5jyz4sAjksmG7/aCMa+XEIU4ctRSpeDCJBl0o1OZCyA/U22fVGBP7eJv9h/iJf4H+I/6p/iN39n/iN2a/T/EeNPZ/xBXXhs/4gLh+hOWD6MeQbuj/AHg923/OIcSzwUf4npOoAxEEnQBiEpH4KlRFxDKMZYwjDQiMBnn1iBtMhdN1r7lsepYA7z/qNeQz6DjEoqMGiuMS5Ot3S3q4rqK3W5ZWFc3A9ViFYywNuX/BKcV/hMAvPbLCl23UEMg4p1EWgF0qJvLEzUI1YKUNX2sVTYLGAqIWrqy48jf6jshbzMCzHIMBrFgMc0hVVaj+0LEtJxcUYK4qP3C0hrqniEKJbdvnuYxbhn1dagsdlX8unP3Kpc5n7BF/csF6sLIOswDSIIpS1G7cFMduztU2xRR4WpbC8VzHPOExVbgxTB2VEGWNZncLghEDu7gGWDh6lPRW8xcWRwQp3UsHgGXHGF/5oS4xBgehDQdhRH8zbDyxR1eMsTdWruJ9GUZZKcG5amFx+5ngPozChV+yWbpviNq/8J/2vLCTWEEAfcDDKGvyBCCAe4B1PUE/CRUDHmBCCMokIqEEFCCYGuoQYkD4GUIOUCBAqEAgJVf0D8c/13Lly5cs7m2D2zYh7EQyf1m3/GiZmbb/AEwG8vAn+0NAHbRBYuKxX1EhJwVEx7+THrX7RiucxjFkSotRaixfgxYijtNIp57ijERQ3KsRte446jtj4HhUuxojl9TZcWF+hFGCgQbAq/mUZSzR/tuGPhJfpIsAehWtfWJqvQn8kv7vsH8wcSnk2VfmVMC3RN8KFU1gJUEKpRkdrxGBx9a10VFSZNAhGdjWrZ6m1Fvb9JQbvETIoeplsb5Exw/DMfGA4gmW43OvGiV9rPOUtNcYqNaotdkS6/BL6aQ5tbTuMKFq4JSFypvmMaNuOYNnuUAKoqiZF03pqIOW/EQMIEIuHCD0lR5aP9yisX/aGhweZYZN81KHZu4xYoBk5gBt5irmR/mc71MAtBxBNNtO7hhxqty98Y2x14FvlnYy7Ll6bwMD0bOLi5bMuIsWFU6CFslQIYLKu46tFz+2aJj1LHAGHIqyA1m3zPIwSmu+CKc+W5k0Q8ylPfbKyaswyrLZ0ELjD53L6T/RLP8AizA1rMMYCEkhIWmsO8Lw8YH4EhhV7lIEqVnEC3UKMCAUsCvghD4Q/A53BIMGbhSDfwPcKg1Lgy61D+laDFD4frlCbJK7X/EDa8FJX/XB/ec6r/niK/eKzQejFzi9Am7W+lNmvajuJ9sVFa3iW7ls9y48xfMvcvm4tsYaRoSm63GqLFqGE8nxLbFuLFiKLEWWSGaRGOZbuZAXAmd+ILifUcF/qWYTnMFvqCMXcVRzB+pnvUR2LyGVQU0DSa4qrGIO7EMGq9zHKtFFujqI70TPCXAgRTpP5oKznN9ItZbrCM2VQXwVKTinUcug6vmJy0UQ7QQpnV/uCB2GWWVdK+IlsCxjMWBeFlFaUrL1HQGBTuQGQ8vUVpbHdnUJSGybq/8AKFN1nzEm0u8WxNod1ANLemOH2b9ku1GaP6iFjSo5vPcwCwTuOFu4OaMuu5obyX5hoFLxFVneqTU1su5nzitRW+8Qo2+kzCw0K8Ea3dX1LLGbN3HDeG3UGGhuuJnJyz7gvpwR1lArETJaviX5dREb6hzipmCiBfJMSIeOrlDbd9SgIKMqJ4dF7hrwdp1Ba5+4ho1UQheXfqN/0MQf83LApgZlfAVAiMwhQlSoEPwlfiCgSsQKgXAgfASvPyQhBzKh1CHuCXV5lgy1XcpFJaVmiUoD6EEO+QIsIRhd1lcvMxTsGhrF8SjZV4QbTfWIbH6wUvD6zhtWU2y1X600i/Cp7mfQeGeN+ZqG9WP1L2y8KP3HA53b+oxmnoCYX27lHNj5YfZE1ieWUwIjpJUqI3BLTUqpUS4Hw7jHMYsWLUaRb7jFv4O47ixseYs3K8RjUyhzHEcQQWRKgILIneYLrECVjVS5Ag5DHcArMkRRY76mR5iLUVs14ilobCIGBT1M1k+pS8RBxbKuErxHx1MzZxLXrTfpLRzkWABWUe6eCDi/rMSo3/MyKx0RtMObxAAFqeCAEUaMMrTi19w71rTUaNm0o7iAFMN1CDgGe/LMqYAH9MrEAriNyDiMcwqlbGVZq3FjbXcGgWX6dwoKPqIbNFnmXElmM+iE1VBpBKNrQUs19THZY9kbxcVkjA89dQYjetpB7A1rzEhhc7iBQ5WEVROheYkF+jMAPQxTGyq3HCKfjiNScBpqXGmKxiLkd0xfMAsL6XUqd2pruZUrPcTQaN3LKOPUCjbeMTG0x/aJpV83LGdOfUCzg9wMmPzN1PpgIreGGjQ+IhMYe5QWX+CD/k5+AQPgYQw18FSoF8QgGpVsCBKeppbAJPo2wZGnBTxaBDEmIFt9xEKH/IRzZq/bRWIfLmkVtwc95qAoNHQYPL9IxnUeXArZT4qWhc7gXxy2imgA4lI1X/ZghBQQdjzui35mN9VmnvLcPbOKl6NY3B4ji/vpaB1IKpaGNe5iou05r8+5m2vdf5Jw6AdtfnxCtIFWInnMahnI6j0XAsppin3cChIq7GGNvs3Myz0agzlv3uf8GF3ECW7jCm2zmeV+ZWkUeXmDUekiB1m8413b+ZdMvzO5/Mx/5o/n+Ydy/cH5fmWrm33AqEdDUBmyR92ZSZ/MIi8r7JTtPuf6RiNlE7R7IA4eyWoZmW6/PBy6V7ljrUep7RixzKHqLFxFjVfJaimY1eYMzUTcMHioKiX8CQXqphzG/EpMxodRJ0RFZgxGHJKcXMkR/wCRBTTKMtfcYVMEVzxLaDVxpm/1EVafuDwxL3llFzKKWrH9ICXDT+oStEJGyis4gYQVX4hdEHGPNwacVuHs43cOm7FRIpAh+SFmaJxcEsYdDBC8hm+pcdUWQzm0FIbr/sShYtnNYgtuF/s6iuML3iW2DRZ6mBbMQviIyFGQa5hSDSJODtPeEUFrxVRFSx74jJy68kduXGJgbXzWogpTXiNhinmoBVnO4j4HOJY2dibgFecFwsy3V5cTYUy5zEEKSsS4pC4qKACHUyL7u08QXSuY0KIMSLzcoFBSueIUga2pDMAXtmFb26lrDAiVlBnmXdQCnfM4wq3iUdCceZ5A6JdyoniVTQAyht1pqK5fs8RIzK0CWI5og0LPiDcBMFVsXZVVKOFveUI0VGNkbal9X/hLhGljcrCNOe2DECMcnNl4PtgMA8il+aGDJnMrFfWUwWENx9lGU7xClH+oIqfxKaoiy48NrvxMFQYUyvN3LqOu8sFZEsBFdUo+o3RWv+ZGF6Nb/wBzB0AtVdWxWDjmKOCvMs8PE28Mb7B9SpQJ81AB2YpJYpa7xGs6HbOEHEaMitXE3SFOyC42PEpDjGrmHMYGzOZSl5dwwLYMZjAXTxcFtqcBKiQAbrVRjExBW5jSgvOMR2J1ncab75gDmFfBEUFLljZRBqEX0scq2eJaNle5f0YxcITNU5qJfUVXqsOdxbZA8weQsyJVBi2Ac2w7jEMtXjEMCM2/DZLyy/MO/wAFikWctQRLTzFsN95hqVPkgtqf93FKA7qUb/iwcTblkXEVY6n7R3Ki3B9xhKzUFnj4LSWHxOGOcc87j5wfUpMsD6npBXEbZccXFPDc2P1L2Uj5wKeohKGKRW6j0F8zPVepzmZrx3EDx2RZSpuI0Btt8YQjN4ceWOkB9QKyQUunHFSkwZ6JfZTaVAGnpgLs/gti2m7fDEVtEMFHMtM4IsZgziEFcF3FdwqUrlIcuoqIAhg8E0iGrdRbWrLu9S4FsBeMQz2odDFwX2dFzmoh00K44jvmTVxhVnExbteKuqiSxWmYW6VzM9sRAWULfEsvQviDDarw4iGGOeYWOKeahjdb1BOhp4xLoULYOonmyvERAF1kYttandxGpo4c5iZpb3q5UGEHeIhVtQis3F4iVw9I8rKmBYpE/FH8S80FDVxol/lBBeMKS7IU1m6jlnYxG0DsWsRGIOShqCSE0pFsVtGHUuNkkpkteLjizAUKcbmV3TxC1BGG6/ZKXFdS7TZ8RN+q/cytKz5hYCy/cSJgcsFWfLiAU5e0FPMFJCqszqDQKPmA2iR4hw3ReoGiQOJfmzRDAqnuUVdqm7XGusXs3KWyucQxApiFVApdwIoGiOBY0xiLbTReDxLd0K5hRNviVyhE7hAcsBqxSZeaxBAtpih5g4UlDSxQzoi48wJ2Lqbq4Nllxjio0l5ZY6YagGxMW9KlE66VmoIXmKyC2bldUmoIEWPMdyt3CW1Wqy1LS3MRgNwHkv3BpUPzmYs1QRiWF3ubmvdwYVVTDM1EI73A/mmBuK9MFz1LRXMSRUqXFpijTmXT5jl1LF5r1DXCvMO6PJBhUHVQ5wPDNkq8kudD3LDH5Y3R+aY7uKXGooyxoiQjd5lmKis4i6jNYP1K9YiFuJpgqUBtvzLJq4XAaijaepw3BdcMVUc3Mq86GOsp+O5QZsY0U41PCVvplF9wrGrBZ9IVNyKPaDff1LVpFj+6MgUx+Yi7C+WUW1b1Bae79y6Gr0zWHI8wMECU1FX0lstFj+ZxiyvKSwtW9qw2A3hxzBbp8DuAoct184iEpTYnFBmNCcDb5Sx0cT7ZjMgFar4YgLpyQxyo5qGQK1zLRklZ4SFlqw3bW4AUm2XVwDjVtSob5apxKHU7WEeiAuNXiOhROumAOZa2pQKjZTH/AFTA0NpGUdfub6vbbTlYmwAq1TMhq1Zd7nkyA/3gEDawtRdsqtcDtgS0bZqCbg3AgRinZLWCdEUGB0O5Wmi6sgYqBuCjqB5osqOgSpWWKCnq2KaTVmOUg6tGDtzvqcr93ghxWruzAQZbgTiV36ZgQHmHWbOnmCGRotVwQIuKmKhhKpWiLtAJ/aGo+64kDj8xR0EEmAgSZM/uYEWzWo4V/wAYEqsuwXZ3FTLYcdQBWWv5mIbfSUp/eYgG+5c4Y1iGAqoQ5PEsOm5bEBNRHTXLBEwZ8xMthmYKpqMQdXfCeWicTYRGliy0xFhVYp5lgjIF1nUBE6A3HR35iUQSzdQAfqVSH63FB2bfLFC6rEcQ/iDRRfcvZbMzXi2BC8YjWTRL2CY3U3GHlZGP4QdszwS06IoDhYk4wRQG8NzhkdZ3B4fiJ5UcFYGSVhwcXDK+JlknMVLYs9ohIvB8KDkn3FJ7RFgOfUpexYM7mFWkYMERLclTJAD5lfT+8zKvsED28w7HxGTYeILv9JZWnhGHEb+obZ+5UtX3KFiJ4YkbcRL6nBOHcT33PCP4TfzKevUctR5o3bKiwSp0qHjH8ZROMxySrlhv9RDEJbxTfpM+4D9odncsvcwhTNdxoNV9RjPJ1LmA81MYqVD9xun1DwGtNy1aWmIRR27g97DM5uYQ1s3xCvRY47lK0Qne2E3VvzuoMehLGIs0CtpjEudFs8nLfQhfJSQWqrNq87iJQcm7YdALZ1d1KLpOXDCv7ROEXghr9CZi4Cg11AorvY/iHkwuQ39cSkghDRAWCsUt9R+vnc5lDBm0s35iMBU0CGpgKy14iRFFYaZfVnILEdg85ilbLrJMgogsofpiTZqjuG9+TGmxGc5ijYVeJcXWzUrArZ4lA2vkgvaq8MXFi45hZWLwVMy1riuJQFG9YzFZpvmpasKG2cu+rwQvPlDFB0ZYWh5lgGlKHMbtzx4gtLqsS6WfuauK2MLxGMsK62eDiGiYe5YaQfPEBxeuSUYoIUuGzUtNpeB+4OtflAIOR5hK7uEtfe5QDnqIacPctA0lYjFl15YFVstvmAMF9JhIVyywpK4gM8PEdRKzlhgU1hYuGG1iiCsEvBDnxAJTS7A3qMFfy4l3F3Zva27muvcAmoMhnUzhkJQBNa7id2FQ0JzuG4u3xGwszjUUU198y9BygGi8ViYc5O5Y4vHiNquPEZiXVU4LlYMPxczjVksGSLV/zEVxMC7pqXBbdRALctbcwUCd1HDgNDL6LwblnMRTER7g6gZiU4q48xwIjHLuJVxLNRtipU3GsYl/+ZmzBVxthZcRYLxxLFOo7qWtRVYauIJ13KFFgR49rHDZPLVy1JiGVk/MHewplX98DhMvmCVKh8oeeIoXmu4vM9yRiWEd5qCpUuS011u6yy5CtdWmoVQwNqTIaw4lIMKywMEufolgrPCMUWLrAlHVvuIsAX3MlZqKvczu6LHVOh/CEAQw/cDGtOoarYZxKFjjKXNtjWW2CulwZEH2y6BcrqPQtI4JhhPcGEF3RYXDrtaaRYXube7F5rWO4SBGHw3G4mtS7bv8xG++jAepmv1Y4InBWoNizDTcl/JHKAVcqypZsG6X5h0ocGUqiPpQBAHDErggVaIimC7tGAtDq8SwKCfuLyK3qBqW8MybMZYYdjVsuiutQGHDjqoikJmxGWvdjIcJQoOuaiDZFSwgXjCXYzOIqlk7lQXJRbEtnMO0q26lZZQ5qXK8+I2DNxgQWnLBvB5mWV1ASA5asiOTEoUxZMhxDH37mBkPYQBlriC5DmptfteCFizXmxym6ghYVAd8QV7+4DcrBM4iRoxK5DO1le2ziDyfQ4ln/stGPVVEAF1mExdwWlUc3B+w8ysvvmVc6t/cx9ssDV+JU8u47pZaUC4Kx42RAovPEECmGItg7/UsCgJ1BxLaiUzYPqXYnIdxnglAYepZ9wD/AG+ozXwqF0dwRASQdvcWIcW8mKFunizZKrFfJiKkcqiKGQP6lEFclwErXTBVVl9xGNVy8wG8U7uNAN9txK9Y3KUrfmMJmaOa4uGedENw3XcpxKGoUhxLbriZV/MpfBLCri5yNQtLyRpXUJlb2wR2YqWxIBQ7hqtM4il1KauIPuKRRcxSmtkXB/UsswNQDiI5Oog6SYMSl3uMcRxKZYAK9xTN1UymF/xLL30mVh+IiytSrGvuVmmArMcxOCuYuSGuIi7AubLtX8SnQLjsLJyTRr8TdC7/ABKuQ+K1FVGJyMxg2FTDC3d4eZunIbplQ5F9/iOvOuzlMAC9jdxHBwC/xHNHbWX6gtDsrSF005tM5XN3bcRQFu74jFPOKwswdBuF0UEwgsbUId7i2uotVQRKQ2bH/qnU2OCY5YKFv3UBC5LcwpFtQj+omlurp+otGCovpz+ZjY2ti/iXtaZou24dkIXIMxnc6eYA2qb1B2zhAl36ZmwJerlms4oajApDrEe7QXYS1TjcAbFsBfDDU39oAUoKqWrfW3uByc808wOeEwrBfMNAcyoo0KjCWWdsuwvGEtAG3DKS8uKjwDD3AjXLwxareXE6FniIyqB+Z+dm/EuwG+WHZuf5jQjR5ViKwo9BKCGq+txRAAvncs8guENytyL4rcWgJlOUfUJh2QizxXi2NVHgoFQ2Ve3fxKFMptok2ItUNid7xKhEoWXMCo/sRH3gnnDQ5zCUgdESkqwjw3jqN1NXDWeIehaWUxHIY8jGYUQFw7gbdm42TH6gVx6iCoBApSrUhUs5+5VU1LmldBm7londykTNQXdBxAo2f3LqDLoNTEIXd3qIARi8XxKb0i4lZaN7fqaAWmjMpsRXeqvrG45W7eXuWRM7tcxGnXiYqqWywU1m8yhZWsD1HAFeVLLhbpWkgjgWspMRpdg5hFMCv8IpSKusQBWDV1DXmr4gpZlqklXqEUXcuau7eCEwcOpUYBjqI1K6zHivxFrmAnENxpNwTB8Yq45e/cu91HdBSCkvniAKsHRK2rqWKuriaotWerMmpeW6ngm0VeolJQ/8hHdRurRFgcEWu7i2pbD32gOTDF5Ydt1WyPBG1iFnGeGKDGa5IimV7lOTHmMVaWE0GAhPRE6cpHLQ9IGWHqMWA9lxpZWxSDdcruItvsRvyHFSwCq3dOSZVHYcxS1Sycxxd8UYjsq5plqDk1kJbKFXFEKrwkHVV04M+03p04zBdVfDZUaoQuKcMpoqXEtiJtZuyPSu23NoAObuMpMmfEQAk5DiC7SuEpmUljFOElvSmBTEKByW7xwsXdvcGwZpV7gg1orJQzqNdystcQQrQV5YqzgvVKCqrg0xZoim3mEr4Yo5m5o8DmBoFcZLhqzXuMaFYiti+GFLsY6uWHKqn6n5CKwWeDUaVvwQAW509kstveBYotKqFSlHq9yyseR3HaU3urjCIHlYYrDnMUjbwKrl3SoX0IQSB4EYBTFXYY/cLZfW19wsNm3X7gJS9mgh6j71F9kMotsSwEbys4anAn2ECkOHASsrbLByEfqDwoGwQ3GiibuFJSZo5jNpatlywKzl2jqhyKyI5ITne44CiixxCKuiXamTqlHqf89YI8mp7bLAPqOKnm+YN8Z3mU3ULCm2CqVCnuoXQZisOSuZQpQ0I6lrKV2JXSg33KEZtmiUMAvhg7FDwShLHFepmnK8dxoFC8MUrGDt/Uzkpum4ipCnmMHLNzM4QVRLnEQlNLl4gHRDGNzFhOTynYQ8ALtKXFwdzLCg8kL2rJ1OFt3BDinmHRQxMhFRoiUu+NS6VTmCg/ghTYbxn9wLlXxHSWDdlShyuW8y1u0aYbWjTmKAlV0Q0EGu3Eo17jtKNYg4rfdw8JfGMQX4ZwIFZpUwGswMaplN5gYS7pgVHK+5Vb8kaMwagZ4DUSNw6QfIsrC1dwm8wNvMSLuaXiJOoZImm0xxGu46rzGSzWzmdpQYUWuAQCw/LBEQFTVjdzKfR1AShuWAPPmKVw5mDjUXXWNyjS3GZ4qYCymCZcq/EMHLdSuDbEoDbmarLuJYl9BETjHkgrgR1dXbj/EQ4DoYkcsAdQso19yxBhtl+YHkctCCG63SRWlFw0bgxScMJg7G16mcKL5q7OI2w20syCUG2UApdtXEKQXWsWl3BXMDqBgO5QSsO3UxF8CwlF3FJAMRyNepYnkJHKc6Y6iCtmcv+olLXnqWVRwYoh3bDg5hZXba5/UxB7DUqamS+qYMJW40IM9IeYGjgh7qjvnM0SDi5kYG8SiqpyVAcEIteADRhvGYSpAt0MwASG6deZTCNBRr9wLWv4QrABuxa/DDaOIDhuNjVfWocl8T0uPFFbu/Ezh4j3AwSKKJpTkGT1F7EMnGJtlQAasgEcGLXAIxIUcnmVpB3TDGUOYdPuGxU7WXD1sRxSWApEbGqjoUp6JUqGUzMYHN3VMMOhFdzUq6boZZGB7lAiUM+YbbV13ARS/mJZMg4uZpxuOoEvT4jsWLGyBN3P8AjuCYNxH2auHj8xMMEvEQxvxDZeoaOJgBZdQy39QW1qGm+ddwgYDJWuSw2ZmagXZMze+alU2ely3UXmoOgZejmVHB1da3BcUo2mZrIuKCXlFMAdxgcjK68Rr1VBcuGYrMLD/EIMKmPM1XXp1HgbIPgqWxNuryRpRLsNI61dLnco71cBG9P3AtOK5hVImbuDao1eJRVFWcyqote7hoFDW4ZHcsUCi5qbigPMRGaRz1GKtR31FzlWBzKTCF+ImY66ipa0S4Jn2RccnfxGbvEFeCHA3G65hmv5gz1cIGdxKWorzNO/hcXKLBq8NRjZgrfcYPbmOljMRUTjXqWrEbZliMqZDcO3VxZgYnDKEJVu4yzcBpjnXEUlrCVIRQC0F8XBu4HMILC2HZM9M8syhoQIK0vEMxu/MVGUF3Al28bmRbAuEwwxT6m0LfVwjaryXGqleYiAQVsYiTcy05iwQ+TLDMoxaVH3VFchqNAP8AuczB9LFLuODWbNEHLCbq10xAYeFmSXY7OluVkThAClzjEU0opqiUl4GWZ2X74n4CIAjB0MMLhrWv1LPTaNlpou7i4JkDkgCyM94iHLI/4l6ih7lOi6zcdYJf3FCgXm4FWWRimLGjykRIGxWFMuJnOsOoUHI4HcJFA0TaRrBsaYkFITVBZf8AEVCSF3TZzL4y9sDAo6ax1CSFGkq/9lupdkaL8sRBAr3qXI8Cx4cykCzYuMO25L7iR3RSzfq/uOk0MUqO2ohTCo4qm0DmPLrSYVn5gGNW0v2EALcgGZcDdYR1BsOG8VAgmGcfcqlbo7hRcjN1LFHDKA1zcoDQtuZYFDPFxI2BbumItDEuMFJqKpbvDC8XL1iutVEqy3WGJgd/xClW6PMEOLvXcGwqitXAFxh7hgfdkb6K3MgrXPmYQFHmXENP8BHJxzPKPLJfwFHXuAqjPUoq5xEoPfEwK4eoWCFVAKOUmAVVfuPjfNQQTSxYu6mCee+eDEcoCl4RLWLqzdnMEuW7GsS45a5PxBZUChrL6gE2DAF6My6U1PIuNp4b1SsAwb7HBiU3zasK8QQApkBuIKk6SS/dVHNHHX3KVNJuJQWocQyKVcsIxx3EwGDuVhjBKgsHjuYLM9xzXfcahOcURVCmLaTULbzB8KtnqNGaHLcW79CYrVU3fcJ3ix3KKIUscEyjgjjNV3DW23UN4rMvnvuBScw57ZRtx2y6WZnkzZhd7mRmG9+IbStbhVYzLzFc3V3B29S4WjogsWlO+4WHUranHyy9ZyMQsYTJxyRLcSxxcNsgnDEyP3BgNZlqodq5tlnYiyxZIxniaE3OY5JegjHurqYDd/mLRdWeFiWqWOMh7hP1JqAS73cQA5eghCT69RCuPDmObYLeEat06siCyeIV5TZWocw1Q6v6gkA0McPMVH7LrMGNRuYUQGHaYEq8DcobiBKgFqLsYYuWKkFYleAwfSCkUOEcwIQS7LMETaKDYKmhUNpn3EAK7DRGo1i8wBKSioLQ33MhRocf2Q6xc3EwUnFXDFSed/iBF4Z/MQXMxRuNhFgtVS4deKqGivlICIVgMJKwjuAMecy3PFF49MFrtUrHPcteFsL4USp1HrURBU2WQfcEqsFkUx1BtFaoDVhaARO7uMiBMYa5mt5opfxD7Q03BY2HfmW6ydEdWuuZaASuYLode5RcWqZJms2QbTs4Zna6/cEdKwwo5vIxTRKdoRNM2vLGLWB1MkzhidlmpR4o5ogirPEptLZipdJ9YgjTm9QMpa5gAEZ7YlBemZ064mznqKUGv7S8jL+8C1wkFXELnCE/7GwRE/vKx27JQjcwq4jJ3D8oHC8etTrS14xFT56nY0gaqCsFu9kGeccSp3uMIcSlEy+3UyNUAvqLqsBxKgwWC0qoFa4ZfeSKyIGA15eWMuohZsOpg4zYKro9ZlvaFKNusQ4NfUOKg8w9uOYeA4FKVNHmXBRasBjKBnWtlZglNV61HZzeqZjKuvuMKtd5xiMCs9i4ArApmpZgaczELLvbMBsSXALVTnZDeAsq+Ym9OeoU2i4UlMyDgy32wKaHb3MzarwypstqYtF9uyCUCJvUpYseP7fEs/xFZTVdwqxqaAjxqFoN+YsmZliFxvlheFbTI3vuYvV9RTMq1eL7il3uYXeGelBAvG5RRAsu0iKUM8wK5fxG9dR6bfEtcFHcZS7gK9y1aPxGiwK2RTuH2QgmTA/qLK1KqpvqBk4c1DKOTUFy5iRp0YhXCSm5fkYQgfsYgFovCXqOWsBL3LZPNcMtLUwvMWsCwHFxUl0SxgubgRljpnZZY29xb2vW4qD3EcbKtVLLrKqscNQa3r/rllKvmAyXeL4iYIouDibzV6qJYXe1we5fDEMnUA0KdwmQQ6I5ivG4wKfUwSCaMwrYQUBHLgT1G/JsZT0Agg3h+I1aAUnPu4ldFcgTl0A65qXsVjjlcDZormuYoqKvLiIGEb4uMq45MxoBViLWNnmZ+i9zGpadMoW6OKhwpaKgbzxHLE7ebiQwCFrBVxUIKtHmPsoeEsoNyplkC0P4jNrIQi6Ym4eeEBtrx3LDHrzPFtOIaN305hACl6g8kw5TMVay/wBQkopxtj+s/MaAB4uLd8rzLpysQqqnUVDrmFhXCwoOblXxiC3F9RhvBvMZuK5jcL7tjVziphuqzuZMTLiIV8xcAm8v+omeCPX3cDJN7MRWBi5k8RtAJYw1A6P1LspbiOpKfEKoWvN7g5P3KJvH8wFHIj8RNXGI2BqLF8CPRdFXglU4RuJJ2nGdR0wKUt23Eq2TC7I2yXWYFDILU0BBVIjYqoDCOwqi+pWSsW7/ANy6fxU0AiBzObEvcrxKdQLgL9xKLQV1iaA3vMBbWvEJQ2GimLjUPF6lDG2F+JiMzS4Z4lQOTb9TLaz9TNcKxmfgNLFCCoyuJShZ7YBWq8dzABXiLXcC+eYrqocX+ojE0rEqM3M8ly74gp6i9xDfE0bzBruYXjMGsNS1qbqXM4Zho5JpTzL2bzAiqMW9TKUK4laDriWhaDaSugX0ykLWIAV1xFFGIZzuVURobY3MmSZWLQ8kEcfcUvDmUxsgrQrFGki01SsuaiFnLFblfmILVHiZufEFStmcQDSowKqOSmLSbzZxHWXL/qjXebNWwkW5vnUzDlT/AMjVWkLJzGBYXgzNdUmmpnD2eYrfhIelYvB5jsvGa0zpBlYii0cNwkIuSupmgdXGLdI0R2y1tUqLzmUiXFSsmRlocHXhhVEHoeYqlaXzqFbuhi5ld5olotkxAtZejzCgFyXHAUfCCd37XARcjispL/Zdw4jHhY6hirv6ioYGxiOXFkrzpWsGyGgutRHN2gyltxiVtC9ylKs4guB9QgSvKyjKhwf5i2aB2PMZDaXJqHCstaoj+g9y6C3xzGWGoBi3vE2RbuVFqvcsZSjCnU1DWDMAwrnuWFPuNKDBUa3/AKihXMKnC9ywARmXgW2tJeAE5eJwF1EAIwNu5xgR3UayBGxkgAKDKvKFAb3XEVQbeWM1XRxDSthMI/KBdJE6yvqVQAjObrMTCm4z+W8EOcs2zoGMspeJVbz1E4gopxBhX1GRdMEuGOILboPmFIkzfUBBjs6uU5EIqH+IoMolQJWta8wpTyw2VuNVw/UsFumiK0FanfuUCjDX1HgYrK3klUOYoMoXqK66qPKncSbAFBuLaDMwEqIaw2TWaOiO7DWCaCUcxMNKqsw0UFusxIFs/wAwCEtHSNoDaO1y44gNOZxmF3FisRBmBtB5iGtFlnQy9haeNkc0Sr7eY4nTOGEihSm6zCTt3Fdrq9y9WVeNxUPEs2wdSgF34jWZsiH1LnMaMVe/UstQosLln5nGXpFlLxA93C6uoo6fcEqNxSkXsViOy99Zgd2VNOJzLX3NO8Viogt39RzmM6lDkql0T3UXLVXiiUUR1n6S1uKzFVeI7t0S9viPaZI8TJyX1U73g2XEsNdTajMpaZd+4vZo4ioF4rJMnIMOCV9wHkcXBIzm8VEioQ8wiBB0RipFpdxQr9YXBKVAck4Y5aDDNcMEWRCmo2lC5qriiUGA+ZSVYyZfuODQAYzbGVxfFxwqAupUHBocQsiipiLRThzwRNasNvMrvVnJupRVwRZc49cRaJq8VDKf7IwDYQXNl+oisvgJbRWtRd2MuLdEvMsYLzzLhLHZZGNeQYgUllTAbXu6lSVu4pty5uUrpOSNiol/cW4G+F1Fbb55YQ8lMFAweTiK5S5iO7WcwBDDq+41cV54gHJ4hlxamLhzMc8oVQ0Mmok6AOCDtGwPcykB2i6Qv6gKjviYBY8S5hVYgyAvcw2cQL0viFBc+JRZzZgJguXD3OtLVxCuLErxFaS/TMBZbl8QNjpdxxBa3FVQyvOoWwA7dEzlFH/YlJbymAGW3rCX1gThiWRdkGvS6MwVGBsiiCDlHjJMjs2x2jDxHrQ4K8QYxHNqWoWQ3Bhj/cpN7jmv5jaGVFwPEvuWy0U31ETw8VCNqV5gkQKK4xqZsKyPMz21yTc5w6gZccxVQo2zHt6hp4lFEysrL9yk7vfLcaGRdb3AzIh1JVtzQX3Hlxk4CLFcPAUalAo+wxCByIw5V0r3LlHAZxAMCvLHohrOYf3glA1Q8zF2WdR5KzSmgibUPOCj8SzbPXcV7K1QykAukxjUbKHJddTA4sx3CYu3Nbi4PL6+5WRAzdLcxGKSqHMxi8NE2HrfmYl2vEvvmNcqx1HbskHDFfNRMdQOP3MljLt3+JljmOt6i5EomdXuU7fcRQqX9QNd+pktf6glu3iCWOOYeHncRvsSzxmHIwe2AyRRrqrbKgGrC8XBVGqUkAW8BL0axzBQMpljp8HEzIN8RvZKAycWdQAClLiV/llOT3ZFEsR46j2Lp4iVrv7lTBxxcazJbwwm6p89QgsV7eZdd3yvqGLumX0bG8fiFZNvFxqaUv8A7MqGbM5iVBQA8Ooll2M1bEtyuxYqVTe5UKpZruAiFDZfERA7qvELeKU7YjZtdlyw8I/mJR04mcWrUSwoNXL5GKN3LvI5igoD3Brh4Sgbt7XEpkt5i3ZXWkHgGiqbmNftDGLL6SytLLywHffcRDEc+ZSBo79ymQp6hsaK6IvK9t1zEjgdPU7eXFSvMjWZQ7HmoASx4QVFgddRaqWsFQKQ8McSstNrRmIpd0aL5l6lE6mcUOYQoCQXJtyektCo6dzEsrAFYTmiWA0Z4hRys40REoazdalRpX8ylQDlaxMEOdsS7fjUvXk8RG9UVhFGDiBVayIZx2zeKu2CBkB1EggxhgbrJKZljMM3GXEbI5c4TUABn45huXHPcN6gFkpBgOW5UpS3RGIU6qI0yeuI6DnDqpgViN+pfY1uuYXFvzC0vR4IaV6jqmEXNQcVV8xbXUHDHgOoFuc9QAYb4iBBc3xuNsF/UcQKb0EuApgSJ1S3nmNpVhkNMdbCFR1RzS3iGsLrgiu6zrqDUB2VOe1ZuYOATctaiMudRH6i1mvEXMAZyQGI1N3qXoHNwMWS4VzEBtV1FaAp2dQlE9DmMAtcdSnCrZY5tpnSO8VE5lo0iq7H/E2QTwGuom75L2RXbB9kCKoPmWURS+I0lscRrOuKGDYK145uHVijhK11EBbBqUlNjacy3YXW4oLdX1Gpj0S7Bd5xCFON3N/XFxlAWsSF7hQtealu8zNn+YutZlW9ngiotVjEpHS+7mDuWJSOLmGL3u5sM1EFONRutg+kQppjcFL0ssbbwx4NB31FWpsnW40OMlwlVeBGEaNy+Ky+YYOGXK12biqurNXELzm4xFy9wstDWCYbmzzHriuMQRuyt6qUFaz+4aFX7RsVan6mDezd5giVtKUHB7h/CJYDBhZAA2rUyxQpwcMI5I2KWeomKlHHKl0DjtBd9CrgqAo9xOUm8SuSEsXSRLUulbJgyNNs/iKqa7rs8SgWwlu4QptyVGKWs5uJPuoO0B2NMDdu2Y5K5HlK8lXmoBbEfeIhXX5jGtByQeIndsAcZXklXd13GNUfUZyioekxJZ6Jy3RL1tAcwFYv6lULbvH8SvTFrnqJqQXedxC7TavUclfq4CEbeyF9FruFyviojbfHBFqcpK82rqU3dDGIKrMdVEA1Th4YXDBbRzCojZzEr5EPcQC6dx7NJxCJ9IXO1mpWxq8QQGG31FsvwIy0uLbAllNmC7alYcuaNS3Rkiy5GPEUCrSFyyjuNdqIrQOJWzDUWxxoiP8AbHkATu5RYKuIDjHfuFd1ZuCCOTLGc3zuLVsxUROw7uXVtSR0AO4ZCEc11AJCk5u7lxbGYw0p7hsOYW37vBFpmmOkWF5inDyHEBEsHiPeqqcP8Qxh4DUxWrBAd1t7jYpKnCRMyvlLg0+4BpAwPMNgCsUY+2LUEa/MACgsK1MNhDT08wEVk8zQ7fMpTIFquoguYhUGRVYsHxMK5pi4iV4YZaArqIvNyRAKCoZV5PO4IQpy8wbFTm2Msuz3EodDo1BK6brVy8lpNlN5lYWeFstUVawCUwsptxDxQuhvKyuLk0PzBLzY9IwoDm2wItR+AcShoR7bYIOLLV7ZcciWnKFAaYKKhMviKrLTlBNheCEro8lywmhrEWMrrBBYFw8D6rMooDHMLOGZ+rjVXUupcUODPMtUVZEom5WYxGojL0Zv3HGjSDLtvxKG/qH+ErMr7j3yw3h5hUWkc0vWyIu1xMYVa3Lwzdbji7g4dniEmdYqiNQap33HSALbYaa8HMtxVMFnEDGZdKPWOYxsch1zLwcDH3LSo31CMWRX3MNFdYyRmi7vjOJd5NVwQUcs5zxA19Z9s6jMZs/tCKIRa8rMwRWnKZi0DIvmhqMu28m4AIAYDsiVXKhqheIpayxbNYzK+acrmqhKauLKj5jODtr3MIZXrY6o8QpZaoGNthTaS6VliNx1UCgY1ccZk5a/MKxRfJwS8pabhrWoYwwbXn3Ef2P7wFNdcwzGA7JYbPrghqFt6ILurWsmG9PDMm67TmAinpG4M7YHNzvqIVnKIVRZzUahnDiogscvEAplZzG0vSBNsxJUV7lG7CvqKMgV+oOpasVYGUwu5zjXMA3qDDOQ+oiOy2RuGB67ggVvmR3YJq5TVo82RZ14TtKdw2g1juoLWVC0uAVTowXpgptGV7eAOoSIwAJLV2bxKA5drCBpA0oQ9ShaWblCahoAreqnKyjocuYkBlqjMqvBlUb6+5RQMvELBdhguJuL1xHDkwsEyz/MWiirYZWDcEM7mDJV7jstuPNalP8Au0RS8UYZ2hv6gBG/eYHOKjGjqWxwQDBcyrKvplOLXeZV0V7iDkMTUS89ygASw8wyAv2ldYKYzxK4V68RW05gAbOJZWW4KLFeYhd0uorar3ccQA/vKSml3AOnh1BrhTiqiYDacxMNWYgKLwMeY0GuXcaWhDGceIBay7zctdEe5dhwUlQpSoOMcxLlgdEJROFnBODV2TJQ5L2qVIrbLfUNRs6SBLaMIZfIcSrVheMXBctlWbfUIXsc2S8Yl4CVGlcGKyjgBAICW9kUr/xHEZHjqMu7fMzc55ixRv1FhMVBqUQFYrDOYd0HcK3tlh69x/NuLaziKwmhpKLVrqL5RZtzXmDaH8sbN5GpmGzjE0r6lgEDD1KgvhlrLPEvoaTcYEtfcfsgUpb8saKlPiNTdh+cRlrJWJ0MhqXXHNKGouYtu3RLro4xiBCjzkhyV7vzMkl1yHMaWqvOYmD7laPwggNnTV/vL4E90qVnaENI1s2jTJKYgtW8sRABsZG/MV6xRjz5JnMtWOHmLXQ4CwH8wmqt1VRu4QKa3J5lK3do8HBEiKDhiiuYlVXOQaihiHLbFL27XxFbgzlu5kVLFZhsmRdVzBWd6xqPgSt0TZFku7aipQyP4luazeqYOim7jTIEz4l4KpyeYpimspzLyFiNYSXDqlPZK2vZiyO4wHDLcMq8sF2p1nMeZhdIlR3AvC/iWOhei5Yw+LmdGBz2zmD3uYiAKK9moGdsag6YxmpVAcFYIO1WB3G1W6hryalI28blxdF6qG5AVT3LW1jgIMF0p3CVMuFy8GrVLtbsWxZTOqqX8GJoTN8SzI84jgZu7m0pTi47kwQqxLSqJccA8QKaxeu5WWjiEwAVThWEWW0SwDVLlmNtgliaGSpkOQ3KgM+42x41BDZtiFzZFomX9RVjF4zmOqArSyNtOpl4i0WNYH+olXljlD1zC2WJVNQ3ZWcSgR58xGq1cA0j37gUICejrELLxjcELGHU1KGtNVFYOheGAwXXRFVZL3ELp5lNdDC0xfDDGlQyrxHfYVAF4A1mFTc0Y7jr74ILFWoWSqbOjqERRvDfcKrYeiVGwc2QCDrDGCN9DUSt1StTEOL2kQGVvV1iNQoppuClQ35jitKbrkjZQF1lNQ03yrzLgLaxa0sRyci8RAA2dcQgC17mIKpxXmX3BTqz9wbGhem+JU1DPcyFirpv9QQBBQvzDJwCAwvDBqqPtkgjQWS4ZKcypwq3dwQ5KY3ANoYIIbviYWu0aDklA4BxxCzkPX94NswHdZlRwkpUteeoa1ZvcwjhiPAjpZwK3nMdjgn4XPEN0j7Nz200hfPiDtaVKGzPLUQ3anScQOOHcVsc2zsH8zApR3cIm1OJnTSOWXmR0kMGrDgkXQFAy+o9LCzvUVc+h4jNkG2LAqBymWFVMBY8kAKsDjqXV/QmYpibilR9GCNpvZfMKwFFMI4MYC3UE2nVYFSyEMo4+5SCrNgY8AStoDGUCHI/DxFtZa1tpVmIqEUVMUOIlmq0inMuBoTjV53uGqz0sncPI0GJQxjGYoDFlTLgh9Rhez6l1DFAs4/8j6wogWg3XNf5ilxePpr/ALE+6eZmsRbQLtsVUyIy7RWrY3W9BlO5QWtL2ktiYNNFZhlLEt4VuVvK6ShBKwH5l/5VQtNeJUjIhzHmAv7m4c19sstbfzLU6eKjTBFgWk9SwEKvDmAwbtLmVrbn7gsB+iCSxU23r6ig4OeJmcrRuLyM3K9YrjuIAN8RwIc88RYpR/InSqwV/LqNKCYxmIW36i8nyg8g+fU0F48wBrGrwQFr+IsKagDl95ml64hIzSYgKN3gIoSPKCJ+sxqFlgNH7ltku+Jea331MBf5gEcluozoq+40RhYrmxiDnlzFo7uHu4P7gzUWuPuLeszAsgkqLDqKvjEP/C0QY44/VxqOI0UQ4JdKKwZ8w28AyjUcsKIFK74llNURrWYO4XPWDUZVNX51O5CN7V26gCRaKgVsq4masuUzJTHMQyuWKtEYiuGLJk/vKmjKahULlM3dy+Cr1cSY2GcR3BacxgvmyoquSmWyDIqeukWJYrXU7W3ZeiURAjynEaua6IkDMyt4IFFj4buOqbaEVC1klYXUJuizV83FYW4pvmCqaXoN+JUReyS0bTOcw9LAYQ3HN1iYdRVrjSL1suTNvkhg+aX/ABEN0bck7QXz4irRavRVRy2WcDL2gNItDfqDUbM3CiIV2QCs3fELIVsisHCaluapz9QOxVq6m0Z8XNThUcg2emZa1RGzvN1lmSot+oKrcaKlFAHOSWLP3LOP5eJYzRfNwSZDwqXf9Fji7/zFAtTzHfkDEstRm9xL5DeWDtyUURCDVmLrUsbWl7QREFq9wbRWVf8AfmKW3miPdN2wiv8AOkq5q11LRQIsrlhVYU03GKhUAqDdZcxQ2cg5IECIXhKIU1qa1g59THVhFlJXIZIgoBw4GWgBRMLEaGpZxHf5GrfcwmUYFFEKrzKrQKVRwidXY5YUDkqsMU1y5L4laLzhsiwDZeBgUifcrKBSilq5nnBVncUnIIKoZWlrCrOQKwIYhsPEvbWcnTFmiwt8AA9ShbqlF7gy9LIH/g3GHCiXpqnHR+4mV6plOPWYhEWrLD1LhdrKLprUFCi0wpHoI5O5YyF1sCY1THfUQpv6i6pp7lqgx5zBKwCLM8VDce4C9g8EQZMvUBTdnjEpFLrcAq3be4Vo49R5r5qo1qD0wBWy79xM2k8kNaOOuJhy57IrtwaWNjV27Yqx1iUXvriYNZnqAs8nc2XkT9zIGLdRx/nUakc3bOuI1xs0PH3ApQLf7iqors1HtlM1Z3G0IKAkdPMC6wnDMF7zURFfVVMDCuyNIuriU6s9xFU4qCeKZdpbEXvMWxX4ZeM67Iqai2vibblgj7f9RE1dcx1bg4iArnPUENU9xeSaLx6lF1PUVjFu7ZZdn1EALXcsK2dJLkNy1m7lGeuoKXpv8wVLR5lU3SdSi9u3dRbHyQvtQNQqBt1MYDRp3NAKIg7NQMFq1LErXSobqq8PqNVvWxjWKwSApQObi0FGi9YIFMPLqUlg3eF6iosi7YTS1a4TEhgdwow1WWJlL4QeWjfGrgYqjdwrsb7xkgotYVuOoAOy+ojnRio3FWnf8zChbRdS1qqUX1CLba3jcBQK6dy2QFbrruYtaIm8kxSVjXUyXkxL7HJxEFKubmItZ+IojKzdy00veWWEV9MUFW7o4jtZbp/ylwab8y62ETmVvRBCmju4dOLvljZzV0QCabhRZrkmojbj7/tKS1PnmC0LaYK1EoVUMvRweGGsme5YNZzWJyAMxWgG6P5llOQ4TMPMcUQVA0wKVLrk5hdKsWY6Vs1oJb3a3eP8wLoK/dRpkRemYKkByVFNNijHOQ2m68TWAQsIJMJ7fLAKIlH1uXAtHH8xT2Tw8TXBlnN+/wARmiGLbVcErUvKcPENy7L2qXJF+HcBVUpQgZEUP0dwSqQ4eC4noFl1shA34yYmQl2C8kYAaqneIxZ4arcuPP6i1Run1cJ6lZ8wwCvbcNDoFcaiCbyWJUcMuYgFuXHEpSbuJNnD3qHsAGyKKM6QzBIA2DjMGNNfKCmH8S1gOW8HB9Ro8KABawdNASv8rFOo5ZzKtbfFvmUlgwWz/szJWnIEqi5QWsaxFKOuVrhMEzQQPECzq9EKIPglRN1g9EwKKL9+JZ0Z73EIcO85iC5HGJbcTbrxLKjvuUqb8R0HL3LpsNF5ZSW5lANI7+NR8MC0XFHXiPIcMtBnMyLHN8QsDOXLMbCO8EHQ3NAHZxMwAMZpzLgzjcZmaFxDovikQ2UYXhjRZFwt1MigpV2RxAHFalG8DOSFRtSX4cvUe3PqVhea/cF+GJ5xGLtLzuLiXRiVeIlmOIlu8Su3/wAiXo4n057gkxq9MqSPqIaDxBtMdMzLZp1KUm6worTepTHIfub6b6hUXdZqEhjF2QYE3LYOXYS1DK8XFVqmBcDzEh6/cVBmqdRVka6jzSw11BLW0buMgGE07ha2VxqUB+a2suRVyVRADKrvuYnTbEi1EvRCw0B6hsF9cynBw9auGq6m/Es1Qwb7mB5aa/iE2b5ogtAKFUNRQTTpbuCp/wAThvNXkj5rFdTc4Yp5ltmLQY9YtplTUAgIzZ3LCGig3HFkBzqXYffUtosGsYlE/AGK7lwzd3upRXHF2P8AiZFWaqJRJZq1xcvIu+UcMAXXXHcFEWjeW4dLG3vBFOzGPtAAvLBhIlacQZHAd7hRR9lzLIqlniWDabrUfBr7rd1HbVhbvzA2KEsPEQDhXlzKgpTmUIbVzcVVS3dcRB5Nr1AsjRyzSC8ialANLuxnIZDMMgAvDfMRGfdygIO6a5lgq1yuOIFeDu4eNy7YyNaxcpsLvrctOKfcul4WoqMINNW8wzlGhVf7j+ldPNVF0jpa1X/yEVzwQV48xBU4tkn4iAOcL/uHtnauYvBQ2gpPv6jrKw0Z12Rkm6nqC7uYHwUcqs5/MYKGUsC32viMidsHcrFFX05NQrYYurfUNebc/iCwJdcfxKHFKr1GMmLuYSvtFwBlk5ZUxRM5jCvJe0uogXjTkDUUq03pIROxuyWq4emKoM+GWuNJA2gx2sabpTkjSqPFMwOhTTX+4ARLkK/qMdyIEVzs9QptnRQmM/uZcseC6fcQa+QW14Of/ZQGEUtjYX1L65RK5+kukEbdOw4y1GCkuoKHV+TmNc0jAW9wMdOqqEMbEzTqEAYdw2bp6JaYw/mKUu6qUJW+u4OSkzhYoVeuqgLz+oUqs3Mwwe0qVM3glVnGYCXdcmpVVFqfRNA08RS22PEKRopBGMuyKGstJZbeDiuIq2xzKAja4jF5b6ghpQPMp4K09RJat5buOtsaxaNim7ODmYFXZTcrdXiKNAqt1zKWi1/dGzz9y1lurzK1/mJ5/M2eI7bjquYgnviIjHRW7l1H4f8AUQB8R2NvxEsuevM8ArcTZvmWVtPnmYAb4xLIKx/EALKfMQqiqxcu1pnmWqTKcMVB11OHOXETyio5RV4grgtKg9rlt4L8RtWccjDAboxUdpXWIU0H4RgHkU9kDExULqApgviC6qg65lgl4vUFLZd8BHAmw54uWSljkTmIhrNZqGGhV0nUyNjziCVMLK3AB/UoBjPZM4qHhxE7gBoqZ9q8VuLYw5MYwN3iAN1brIxOh9ZNbxFvAblQta9Zm4KlKNPlhWNVO61GFaLp71BklBQXa5uNnXnvmNRwCvOLtgcjuApEYYsL8jCKoNIPUTVC51y8y6YBw3UdaI2mPuX1ayhDiWW8rlFLq2rvEaBu1/E5VeioTXhMg5uKTQPLAx31xyQeU3xBvU5gEFGthq5dEoWtalFRa7Lfs4ikorRXcCssu+PEKhqy6aiKDOlXFTX1ZqCCuzdBqLF09aMe8pedsClJ1fEoDvQwZCq3/wCRZgy7VzKjTQUku2UUre4KCm2BAGG3LHYm2MxhL6K2LBV74u71LBB1YsfLHXulmHyQCxY222hqBgbK2SrHHYxLW8CrRL9TAwE108S97W5gNMsvkPuKhoHBuvPWuJZl04QoBJVJ17gtsHNFuYxFKZoNRkWqrHk6h3WoNnUUth2bPzNmx8jTmK5Kqvyxih5pgAabLc5rXw8RKujeLIbVvPKCcg4w3Dkp0xcysBVS2SypaM5eYBREeWplbH6gEqxd4jdBvBqoKs4ljsXV+oxgDNpKykKAjqq/Urh7dBPjmZsCRYHPqILylepeCXU6comf/IKGKUjQjkoz5iFQWEisb5UZg8dX4KrFcn/MsIRNFVFrTeWyO0DdbSoG9+AlStfcRS7fJB05u+9wtnOyYs5K3Wput1eKgVV3kzO7XozcvWX6jq2zqF2yL5lIGvURd+Gom3l9wNxR5K3ChME+4gZvxLbC14Ymzm93ULZwB3G4jx/MumMjvErbd13GvTdk7Fq7hitRyZyMEBAHjcTI1paylHaReM/iUN9QAN0+dxAZu/MxMfXmBT34lxeJdtPEN/SJot9TrmN2zUD/AFEvHoZp21cRCzWmLvm+Yy3XXmIVjAAwXQOoDluLQUE1XJOYqJg6nVp5IZ3dJzNilt2Rm8I4lC1x3Clxx4hp2aczVzVGJlCWCWxg96gyDld+pZX0XmWljYcbiCG3OXUUKY5OJYUnkzxDdXF1Cou/K+YwW24IzZbjHnxHW4NcFtsYcuTEWoAY3FV2vRLCtAX3mYjTWC63FsGKcXmUBd+MjA810qHkve+JXQQlemriE1FFkcN6hLZHCGBQZKu6iJcw5Rnt2rYYlJZdA1SpWDYihO0qgC/D4lDjGP0DzVw8GgTIWmMA4YumMS4GbWscQbcLWYhRTwZ03KoRu2ZJkWI4MZ4lEzYcMwzXytgq8xsoq4gAKEC3UFWAzaoCFQcA8zOFnl6I3ojbxj8wSlA4qXMBNjvuAxgDVQK2xd42RKqo22aYZroK1rcubUUGjZBG2ui4Y7HG8agmS7Y6MIqHqrbvcDPkKfmoKBu2dwklHC83EQtriClSjB0S06duY1btb+pXBbz3DOC+csy+hy33FhXHEtcPd9QsBpuzxHVjbfqXgYXkIEMCvUNKwaplIWKyjDSgmrWgembDK0ihtqL+0J5CabYFBSnA4ZkFJVhggFHG37hVzFbdsGUyobyoUWbKqKgZ6KXDBaIX9uPqGS3bZiNkSjyf5isWm2Gu4CmkZHYzNQClznBODcScc3rqMLxbsvUqhatN3wzAFAbtjYEOd3mBjocVqIpwHHEawbzlgKyUZBHMFfsCUHCrvmNrCmMnU2CXScku8iPmAt+CXDB4lots5uNkdnIQLRBxmMrh2OqHmV561bs7U9S6HeSpKluR7x1BrGoIlOP7Yh5ujQutIdwbmBa4QgPOSZuIOXME45cu4tgSh+YaCYQ1Eoqje4za/JG1AyC5aNJlZfe4VT9uIgpKp3nmCG8/qChBVl3MVcbuaGhPEyH2YniYXc1UY8SpSXVamwu/UdQrjmKGHRuCLiw5uUwNHDGm/wCYtU/cDj3F53jkIWQUEIwuO5bXN9y4Ry7GdN9RW2OU0Rw3k4heRjMq1vcoox9xzcRPEQIH3E0EdwJuD/qJmplJ+aLUZdEeGDwiYthxLGzCcdzdMLrqHkV6quoA0m8QoKhn7gXe+ElOi1jPEHkmDvNxSzmIAm3XqUkoPqCkbJUNmebgyBY8RFvPiPEcmnY+YxbOP1Hy9IzWBu5cAYVg2ZeZhYRfuCIGFWjTGAj2dR5gDDLbGqM5i7uUFf3jVGhRHiMYHDWNwhUpMCr8vmcciM4Y55Cfcfiqw5DB7dfceFqKl9ACxjkmpGrq4q44DruE+famyEgzS3unEzHefKOnWsrcaWLcbBYMuxbWJT7IOKZ95iqrBqqsL1fphEiaqhWrG6ctlxIroOQhWd2onmCOolSwsrZVY5hzRcO3Tda5D+ZghBEzcA9j7IUHDDV/UG6hNtmjcvGQehWodEN2O84r6gBLKyGbiGN3dX12Q6q1t3mLGDaPL3OhgCiShIBt9Kl+tGgYjoGKirZus3DAvohVN0gzf/YhKjS9NTkR/bFWC/gJlLOm9wmWnCVVTB5bWLlvIrat5lCCgq2niN0YvwQuWs9K/wCIJBNveItDG3J56hgLXBhEKLvxEGXWRlo5qujc0rQw3hnJWB1UqWlFmMQK03q651HO4rCwBtqE1zGq2g4oi3djyBlgtUyDKz0dP94DYLpqaPD+UAhByC9wZy1vcE0C2npiu0OVhV8XxFK1dJvwKwUUKmU/xAXlog1iXArbd46mVWtLEWsb+ogK2DFKh7aiIKbMu4NwACl3cKCpaxUEEoGE5dRW2EUAGYqopQ3VRJxdF1AqRKx6lg5G+cYjcUZVUu66dEvdWi7P8R6CK8yktYuqvmImlJ52kVhXZjRMGDh+Y2lMcZTEVQrOZzuiahd2dVUEhFeZxXVl3eIoUtANVuJOL5jmOYOobVBGqvkTPHcrAWNaCC08CvzDx0fstMSxzJZVKyHVkqkMgNvEOangOo/MOMylEK2vATMAps69x3Z3cSW1jnmF7FrdQx/KUq0dLFBkaSKCslcKjgrM15ahVGNSoZaxkjiOQeoigFXiJZ59QQB5i3Wpi0dyqNHKZtXnuKvHfmZKcuYUNb1MDz5g1as7ZYaZ6Ypc/UsNUw7WYMfMwnnq5SO68kMtFNauKjB4lMzBG4u4mFbgcxtt/UHMfEL/AMWiY8DHusbiFQibydQu8Wz9QVHDEMVX/eEsXeo5NmCeQtM0xOlTlhRZKvNS1VZ8GZ5mR5lBsoXNS2Db3KBoniPCRavEGAnKgjCoS3F4gm8OGtOf5zN+6WRRAavUKK7TtFsAsyxI4+/7QzLxRwk8sCMwHsMJarWuGEbJhHNxwRVaifi9uYDZtm2F5FA8TCjfXqGrWy6xG+fUPam6frMDuyoLsCHea57nDDCUNV6u836jFeLcOQGkktAXIBRQEOarNykSuVLBBTTu+YrLcy10FZ9EylHLgGIlhIEbPsb2Q5KycwmQ8Fscroe4xUcswiNrLlYbtV6I6IHooLBj14xCQKXLiSv2xuIyJD2FeoKSXUAxjv8AUMGEMDBzmX5WGkzCuYJlupZlI+zzBWzrCogoCPioZDc8v1FJvLo1RBtury9TeMllWVhjBQZ0o8lzLK2xWRrPJKUjejC0yRNaF2xCKnW7IQ5sOTuKI5Xg4i82pdviLQ26qD3K+YqtyHUfIapqupZWqKgxcUJExa8zIJigqwzf8xFDxqcHL+ZVEeDnqVAGuriBYC/zBQyduIG/LTBVCBeCBQFi7Uls1DuDXGtqFEcgqr1VQbEBa3RG4vtxNoprNovQX8xQTRtsxEIZLWJmoTa4YTKleSks6bLmErBMuwGHYEAXQcOM19xVpG1YgrqIKx/8m0qAUM4eLipVkZv+8PfsGuXL6GX1KnQxQblTCtmZKptrhG3B6R/iExt7NzWZb0u5wAWN84goiFbcZlBZZOQBKmhoZx5gKlrYUXULTYLsgqjp5HEQl2+G+IOSL2xMAoGcrz3KypqqxuWRRfPBUtipQzIq29FiLMXVEc7fdcSgO+ajQC0YgFiODuZPAW0UAPNfmJgbYmEUaFjZe4fMC5hg257T9SlLCKc5vLBQTB0t0vH3AHq2zZ4zA6SoBzf/AH9pc2BVbeJdVHGPM2Q+HcVciuHjsP0xyHPluMAhZ5dTFG7KhpY+FhbuvGYWDGeZkAmDtpN9Qio5/iWhuIBDfUt5rUpheo1Vrr1EZ78zyeoltOswtt/7LalyywcxTFtwDA8RD5O4OCtRrvEcA6YhZ3L2eX9Sw3zzMGzVTKhuoAPPUr9oI2usxOKnM/V4IhBustTG288Qu71cHPTCjVXHEftsjT/yXGxqMQMnepTmMqTN8x0NQUhxnETd247gs5PMQjqnNm5RJWWpXVKpo9SucjDcr9WjrxHitQ9y1Frf/XLRcrggGFrqmGCgHLKUw8juKJYLvlBaovJNJzZKVcWcVmHNJVKriAGC7C9QTNx3cplBsuf2qGUNXuo1iN5XQUYzjvVSkke5uuAXVc1MSLUtYJhz5g4SqK6sii7SznxEhRWFtGq/hjqPg5XiBJqHJL65mkm1UtpS1to8nH1Gv4UqzR14wR1a5cdjTiKPpzuU4193BU1FWim7XH+5fmoFLtsK/wATCc2gldVuZ0zrovAmI0VXkHMoCiPHP5iMpAwLiMGBA4ZiTFUxsUNC/NxDQDCtm/EvFAY/Fepj2iSrOVN14mQUBYL/ANrziXOW4UVXvH5gOhKv7cRARcuvNxKTd80zBusVjmpmmlfIXKUIBbfMLUZLrUrfkOOkBU4VLj6mMyOKOYEQUmKRuVrimwbWIcrTJx48x5A3I06h6QSvO+JcWIUEQtVtIFFIgUc3CYXRxqUEMtyN1LaDdK8PnxCVKmDT+4LxWOFEUG1wwH1Ly4OENMp9gNbzEQLltNePEcVbHRAP5NL4XxMohLVkXgvuGgBbVsHcEiHIVWSByrWSLkEUNuPcqDlopiVT6AG339TMxZC7v6hdOII0HiV2N3XBEz6lqFXjErhkthaIIpYpcuUWd6U0YhF3DjnPcQ3dNWbYdWW5XqI4SrtxvmIBS4QRgClEu/CWCCONS5KF3TzCX5mHmLxNKvBqXK1TAdxZEQOo0oDpeGCUisMpFckwNUTPIS9alY3b+pTDh3iCZUskugFxAClvqWC7r+WLyHhZd+z2Wy3xxiXcLNzzJKclb3th/gXOW7sBzll8QvLK5oJpMGL3WpgUy6mdUQkWuULZrmV9a37CIAqMNbp2fiILpsDMKdMAQF52Z8PEN3J7TiFgs9DMMhaXiWq8OGPYv2cRgaPq4gH1FG1s8RVFKh+ItWDXJLv/AGK4WxlQufqGzl7hgYy5ruIsGL7lhOce5cc5fMQOliIscOIwGzxFaMy468RawyRSWFRHHUvTxPyl43qGeoi8M0btYJTj7l0OdwLdKkxVfxKPv9wP+7RDl7jgFVzdzNUEsVh8QWcVCjKW4IW5/UF+o1y8QBs+pa8ECkZOcRbv1LnbhzEWQGKlBeSpvPOYg0SMinAY2zg+FJklaIUGQu8VZAkruEm5mbZtgpUNDfY2+2BSG6KaKzMo9iaiKjlc5haQ2ZSiis0HKxzKvLc4phql1DIaTGf5iChVua4lKaDDV1Loj8LfmVyEBVNHmUo5vP8AMEpqaMo6SBomuGKFBt0lAdRC5i3VQwEy5VA12OjUXUUC/olLMv6TPWSqyX1cuKxi6xCCNnTuUsywAOuMbjY00YWeWooBOBco6dWD3xAuSLKy197lIZzh7DarlmtvCu6iAV7LcI2gGu5TmPJBLs8zMab7Df8AeUISpoLxqOXRcIdn3xCoi3DePFufuMpE5EsY9MfFR+8ACBs8+ZRyrPljsNNC5eBDuJr5eOYhF4K+0EW+MdEFQSxw5gMLLPqpQ6ULjtCOStfcbCWA3uMui5GK+9Tk5ECyDvO+IEmBvagVvepeWRCmBjTzmAosDZoviOKrRSdZqYSXren/ABDA2Ivij3F7bIk76CDS220a7YASE47Cv9xa1Llef4gYsLFYD9RK3ENpqteYueo0FAKAlwmIarIW9o4I+wWwWldkv7V0bLn1CBWrBtuIopAFNGJjUFzeISpRFu68kulU28X/AHuNs95Q4r2wfmnbR4iICDY0eipXEAYqU1hyt5hSuLaa34igZc5agsTVZrUuvYoPdSwvLwVcStVU9MBNmGipYKt3jFTIAvVhcCOuZwiQk5dVmNtLKsHdxBLCjmOFZ9nEqlrHNymsLfmIZyWVnFaGz8wiwq9ri2IY4HcWmUiqkTW1Isi5HLEFZebip/RAKqpxe4oN2crqJ1Rw1sdkrjrjw2FjsXHEsOB10pDlM6uYxOFN42Dwd+o2vDsKt9wy8V6bf+JdVLAXbd6gxiie16D7m9YcDClXDZNxTniU3IDX/MdgFd3GFKwtCUe1jOyXtjn/AGl9Xrt4j4NI7jyAqoUG3nuAOxl+1muoF2DZ1BDWzxAC1B4NTMpolgB0bYmg3m8SqAnlN3MdVg5i7OyYMZl15l6GotHmaDuHTcxwgK5jkUznzDIgzTUzQTUrUcG45hlpyzy/9RKGRp1zwLqZjSuoqrDhV2wNpmvJLTiqg28xYzV+ZdJ/LEGXzKB5d3qCl5JapeJlB/MTIxXPcLticV9niK0FO98ywNCmuvEXnFt7uUotXL5qAsJQ0FktAGL0m5DfFSpBw2BcpqmWUVM1hNy0W5gLvPCqhWOxz5YCyJ4FeqgVDldg/qZW7CqhRanY4jGQwYWriijD7gCrweC5dsrig4m9ZUt7Ya04pzMGys7XUQBF4OWC5RVtiwgxsN+V/qIrClMXNEKxd8wySG2+WPYAZymqhFt3g4oz7ZnKNmS1jnxGCFGIo93vxGwPEqjqo4Cl6TTFlkBVAfr/ABAcHKqO/UYqs7rcWADiiICiDNnMrItrasZsTatD4hAb+i9QbjaTeDPFRxlrjF4ioe73EU05LCISxdW8TA3UgX5n5Dqqg8xPpHAt0URAFUXit3LUthjiQq91A1gDtmBtFwaWIC2FPcHYW5K3M/YqhtSrY0dEHrlgdGwoBZxV7piZi8L8kAsxim8b/wAwpusMBf4q4TtpdXWKuVAOLF5gRavN8FcBGNrha0t8LxCRfiLHuYS+FCYfxCBkF0DTWqwEYPBBAf5gigwYLc8cRFhkNrp1GcWyF6+4YroXFMd3CAlmhYz28xGWWpUWU7SEtk22Z7aiLxQtwVHtVgdFN/WJQhQBZzrMIuQsLT1EIgVaODOalm4fHEtKtcDWo00PJECPRpOmQ637lxCnIzANduCrGK6v8GYZzILBMLsqIIpG6cSyAppTLLoBhv8A1BirN1c3WOlt1UGAFaxljsWW8u5SzInKkeSF81xFeWeitzmLlycRJBmzNkYHwuewesQdni+I5uL+40RoS9EvwB5zA7gWWyWgA8BE8rcoaWgcHP8AaKAhlyNqAF5rMAB6FAAAefO4vZcGNQRI2n2ajqgrhjHqYnZYUstuFxzdYW2v71LJxG736mWPLVoCLNrTYDiChnzLtfDBIFjZevEdC7DETajVaxczeC6O4Cja1uPSi8jDxKJlgZ1cToOsSyq/uZTeLu42vQzhmpQeN6lWJXHEbNPOoVWsS8JGmjUFcS2WpnGJbxDCrlZdSqDZFxFvzCj7lhcEaZmi1Chu76Y3af6iFu43zBA1mCt9zCJSLTqZ5HnuZG8sLplFAldCx9ywrDdNBfUd9fmCv3C6rbFYnMYpZgIemS+4Vpw7lBQw9cQFA1vl4jpma0nMK4tGsRwNU8xQgzzca0w3TevpjblAMFamznHEAOLMxEANV6jpFVlxzKDoMV4lJUQCgoq5dBkuXrxBHA9o0KNfcVrAYuWmK9qaj0Gd8sDL6adxCtL48QzEsZVMMFurlTi1F3cOxKhgeY1yHdszUAea1FalF0NRQpM8KT7gDVvTuAKKvLUzRGC8PhjG8tn9QhAIMxRy5+n7gJCTaXuCmy76xLlfSrc8YqFdt2PMdAZWOQaPRHBBxysajiNEx4pVBHaKXV8QCC3No3uUwsF05YjRS3BGDtihVoe+SDYaYwXMAGBb8/8AVFzbeS7hlQPUa1eQwOYmalq7e5lBtzDJizEEDLLeUUUgHBgbz+ZRRQwHBAQQwHUvsMO+GaNxhtPOK1GZklqmDHHcMWgtFfrHjmIYhVOABvNZgsuYDur0OJT8DgZhHedTLYQhyd4lAGweVXClqLA8CnPc2RNUgdd7qUoC10Hq+ZeNWsIjVboMQ/s72givhBqloG5Y0FjZzcfVutA1Wed3LQEHCLz1uAXI2uR6xEN+qBwM7zvGvMxnDa7N52SxVCuwN9S6rQG7bt3ZfslyYAt1434lgVVBKoNwIbW1Deq/3Cbvkay2yii4u+X4lQ3ZwA/v+YqnC2WNy5KAzd1eY6Ftfsgha7Mt8kO5G2/5iJahyH3KCKMKtYLRweTicG0yoR6VsVxllmAtMLFXuzMXI2NWcSyY1aSWSYy8riHEfZG7NCbvVSnD4XxNoq1xcXJ4dzPlXF9y7N1zmXYu+0Sy99xqwUzHsWc4hin8xFUGM3n3HtqtUpVUz5uRynmWiU2sLuij1+5jqigDH9AWvqAlcrb/AJmdhAKgzqZQJp4ro+sxsgKVi9q/Bn7iUxSVwg4RDKCXAfMU9nOSDWhbyAFWiyv5i8pcoMCIP7wF0xqxg4Cszqn2WQQWodl0MKGIgVxRzEqXRcotXMRfBySwBWDrmIzdf4ipisR/HmpRNzGosdxx/mHTnqLZPQmpQOuI0bOsx7qWLOCtx9QaNfmYXGIgMYmRUEpm4/8AkT+x80y4vqbzycQ0l43FGT9S8nnxAwKDWINNRKIOO5glZZgLq4PiEQDWNw6VFaOeoIstGWEc4mdGiFLmvCELGl73EyyZW26NMtrhNpxHJl60wuGN3WGYFRm4dkKNlGdwoZEvDDQbaCjFQoVoaf2Sqhe7tnFANFsaadHUEBEF24c+4BQWvtUrK6TsYN0NKw8xKCcc4qDZ0NYhhEN6SyItwW6TgioIHPllC1ptYEuhnJphdsDWzmWgyGaai0yBoyVembEQ4UbIECzJXleLgoAguUEwV3uA2+PLTAGwrhNyhErmNcFDbzKnSag89SkbcVmXArjCBFLSU95g1WQziZoUGlTAUfAUxmMata73X6lwS1MaKC2YmcyU7lwabwVEIvRdrCqUvEQ4DxB8kduSW2fp1C3WmOGItId5i+johZnPMuq4oGn6xC+K7eBn83iXXgbi6Iq1F1vv8IMV8AGju7JlEdYrX1BSSolKXy8wBi1KALfXEeu6FUf/ALBLsp2D7O4vUUIqBV8yrtaSQ8XxCVUWcn3Fk2QFfWYsqgYR3jqax8MqPK4CioHt4/UAMUrmFe7mKvI3a+HgjgcFLeKvzqIRYAlkHcSGF6GuqDBGYODJj3q/qK12y22sdfzLpE001Xfuqjozu7Gi2r8ywCoqEHMHRcPcJDHbkP8AqlQQXZrgMzAleHFwDwASiNQpybtZolnY3pisEAc3vuLYeFNU1MM15UzcshODlLU0EI/73CyrjCQXhU3sIpCYO+4qiRV5OoovU4OWUix5rEsqVrdeJZsJS/TASbsbjF5SNOcS4nCvmKYq7MZjaYfoajCgD6l3gVrMLK1jVSl0pnN1LLjPCE0par9xZyIttGpbEVyMfQoIuaKdwm9CkLpx6vjzECBmoIkBgePTAsw1jJeejX7jbQg3kcIPv9QTWMxRbDwP7yiSEDlkqcGNvUTalbjiC/HMzKkGBlNY/n6liwKOHefzLFq96sqK5BMx9QqE4UCsbgL1Va/xKV1Kuswh2s8Rp3e+CACjRuLmyliSvMSg0VKlssqMUglUdxoo2v6hZ6DUOwLXMvFEy4ijVk2JgVq5l5gsBlK2zhuOi9RbfuebvEKuNRzTmYEMLnxH8pb/ALtHxPq0NOYtbzA1W4gqBDuzxAysmRV7YFdYqFOH5jRMXaoYPUMwsPMur28x2PUpoNOYIrZqNFDHVKMbhaPay6BblJqR06Yje6x3FhQSdsm4jROtI0MrtpKlkrnKLLOkudDhjjXHMAZ+EDTebhooBaSK7lvfMXDeMRm6njMzUrevEwXA3LzfhDBRXnMXUMFjBNjRSvUFbVLmpbxPDC1reazEAgUUHEBmgqkTcwAudOIQsAhUtIN7KviOxmCc6wX1mGyARWALoPcK6NQtxn/UFp87ipnXNVcE7ZC9y8TBXEuta5JVEOuYRzWpXuW8SWGEaEVd5LYf+7gTPIU40YRwNSZgJ1mWXJuVyaSyLUNZDM27bp7hHytyXxBY2ZzMkBVuGGJt28yotG5V3HBMllJA7BuKMMS/jFVQAjDQGKjfmWsBNoX2pl9YllfsIwDd0eYdluapjXEo74DQfy6mR8OlX1FPYodcyjAgAsqsePczhjg1/wBiJgIyOWZxV1C2F7/tBJWSDOba1EFIg0KXwL+4Y0spVhV56zqMcsau3ZV1+4N8bMgJrxrMQL0wU6/Up/x2RYP1LKJFh+JR5tAOW2v8wMdFFZnU7C4IXzABbUBT3xBE62FYviIlUErJjbGy3xxAssLFrqLtS+UQFCNCwCXFLu8wBAIBYvDP1coHXldeIkBRpby4lDEW1uWuokQBW75My0nRoDzGS4OKOHMC5KKUrqEIEbDqKkDVuMaZdi1ebTmVLlqtVAKh1cWA49ZhApxVzHDl4rEspiwa3uUNDblI6pi2odu4KheGsSiFVWZojyPMS2UB1MrD8mVBluIeBngzLNSJegcXxDlJcYRgPxxA9XPalgH0EvKXdwqVrjbdzGaSmAuhZ/fLA50RgN5A7PxGKWAt/gVJzKDDNjeALXZOBITYK6+/1OmxMGU8ysaM4NZ1iYyCKOx4goghtti2M1uNZvBOi6xCAihZlw0ubyxItxXU0c5f9NBL0c3uKBcEEGNYi0FZMXPHURRTUq0e44Fi4cagvXuYIQWeNy17g8PuDHn4FZC2RzGwlmYqrzG/4tE//9k=" }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOy9WdBkx3Um9p3Me6vqX3pvoIHGvhAECYIECVISKVHUKEae0Uj2zHjscEwoHGG/+sXhebDDj37zo18d9oQdtl7sB42lmdAwRpJJiTRHBBeQ2EgsJNAAel/+tbZ7b+bxwzknM2/9fzeaFLvQBOsAf1fVXfNm5jn5nfXS//g//JP/+gvPP/ov6tpvYEUrWtGKFqjr4uSF773zP1VfeP7Rf/G7X3ny4Q+7QSta0YruWjrlHP4bt0IUK1rRij6I6rpadwB92O1Y0YpWdNcTobIvK1rRilZ0KxJhwR9yK1a0ohXd9eRWgmJFK1rR7ZD7sBuwohWt6JeDVsJiRSta0W3RSlisaEUrui2qxBOy8oasaEUruhXRClmsaEUruj1aCYsVrWhFt0UrYbGiFa3otmglLFa0ohXdFq0iOFe0ohV9MPHKG7KiFa3otsit1JAVrWhFt0crYbGiFa3otmglLFa0ohXdFq2ExYpWtKLbopWwWNGKVnRbtBIWK1rRim6LVmX1VrSiFd0WfejIIs73MDv/OmLb9bYzM7qdS5i++yq6yeTAvrB/Vfbt7y5ckREmNzB991W0O1t3uPUAc7yNY7j3+Xe4G5j5g6/DjG7nIuaX38MHH3ob17udljHfVl8snPULu/+K7jxVzPjACfWLJQbHDt31dzF75yXMLr4N7lqsf/Y/xuZjH5Mj2gnGr/4lJm//GGCGO/4kTv3uPwMB4DDH9Edfw/itV8AxgNbP4vR/8Ecg5wDuMH3jG9h//fvgrgMNT+Lk7/0X8IP652tqDHIPXwO0iL4YzfsvYvelb+Pob/0RBkePLuyOiPN9tFfPob1+Ht3eFuJ8Arga1bH7sfHMl+FHo4N9EzoABPIei4iPQ4Pxi/8GzbTCid/6j0C9NjG4mWB+8XXM3v4hmq2rgBvh5D/4r1CNqv5xXYNu+yKaq++i27mCMNkDIsOtHcPosS9gdPaQ18hwAIdb9MWFl7D7g2/i6Jf+CIPjx2/7efa//2do5yOc+M0/XHieFd1NxJzUkGXcjBH3r2F+/jXM3v0Ruv0doBrBD9cRuh34oby+JE6vY/fb/wrN1jYGZz+O9tIbMokY4HYPuy/8K8yvXMbg/qfQXXsTTCTR6u0E+y/+a0zfP4f6zJMI2+fAP290KjOaCy9j/OMX0I33MPr47+LIxz/Te5bm3e9g98W/BrMDIoGZQUSIzQTNxR9j9u5raK5fACID1QBuuCECrdnH7Nz3QRv34cjTz+ZrdjNMXv8Gpud+DEaNY1/65xgcP9bbv//9P8P0/bfhjj2Wt4cW3Y33MHv3Zcwu/BTcNnBrJ+DqChEjUO1l5eaIbus9zM69jPnFnyLOZwA5uNEmqKoBMNqrP0W7N8Hw/v88ywNmNJd/jPGP/j263R0MP/bbOPrJ58vOQnP+h9j57l+AA8CRtL1TTF7/JqbnfgTGEMd+65/3BCp3U+x/788wPf8O/IknUr+uBMbdS0sTFvP3X8Pe9/4tOAb4o/dh49lfx+iBpzD98Vcxmc5RnzyF+XsvYf+1v0GYttj83D8Gb72CJhDWP/EbaK+8jvErf4N2dwfrz/5DuO4imouMjU9/EeHGOYxf/Tqa61ex9vTvoh5MsHv5Lax96jfAk8sYv/0+Ro9+Fn44uI2WMqZvfR17r7wAqkbgrkEY7xS7I+Y/+SZ2X/5bQT3HHkF9bBNx7yL2X/sW2hsXEGdToFrD8MFPY3j2KdQnz8AN1gAizN/6OnZf/i6qY6fT/cLkBva+82dorl8F1QNwO0Ns5vmW7T52v/P/YH7pPABg+OAnQABmb38T4x//AGE6BqhCfeZJrD3yLAYnT2Dra/87quMPg7p9TN9+EbPzb6DbvQ4woTr1CNY+/nEMzzwCt7YJ8hV4cgU3/t8/hjt6b75vaBWpfRfkhuBwSF+cewG7P/gGOEbQ5oMYnDiKsH8Bu9/+12h3dvR5dhGbJp/W7GP3hT/B/MpFeZ4H9HneeQHtzGHz6c+vhMZdSNXSjJtUYfjo8xg9/CzqE6dBBHA3QXP5PaAeYvdv/iW6/T1QvY6jv/GfoV5rcP17bwD1OiYv/okwhKux+fn/BKOTa7jxl18FfI3Zj/8dxuNdgDzWP/2H2HjoAdz4i38JkEdz7luYvrIFuAH8qSfgh6c/uJ0gcDPH8KHnUY06jN94BaNHPgVAVvfxS1/F5J3XQfUI3M6w9thn0V54Bbvf/3eIbYA/fhabn3weowefgqt878pxchX7r78If/IJDI5vYHbuB5i9+wqaa+cBdlh/5vfQnf82unAPBqfuARgIexex+8Kfot0fC1NjgNEDj2L88p9j/NYrcJv3YuNTX8Lo4U8mtaa9/ArCrIGfXsb1r/7Poj4MNjF64ktYf/w5VJtHeu1iZkxe+zpiR9j82GfRXX8Hs/dew/z91xHbBv7kk1i77wT2X/sO1h75tJwT5pi8+hcYv/UqqB4BcYa1xz6H9tJr0hfBYf3Tv4/2nW8grJ3B4OQpMANx9wJ2XvhTdOOJPA+NMDz7MMYv/RuMf/Ia6rPPYWVwvztpad6Q0YNPY/Tg071tYftddNM5gDlidRqbz30Fw7OPw4/W0V56SQ5qp6AjD2HjY7+N4X2Pwm8cRdj+CWKMADdAdQobn/p1DO57HNWR4+DJJTGWMoMxwPonfgfDB55GdeTYbT/n+jO/D+7G2Pqr/xX+5BMYnjyJsHMeey9+Fc2NGxg+9kV4XMfk7Tcxf+/bGN84D7dxBse++A8xOHlG1I0DxJi/90PEpgXtX8CNv/hfxK6ydhyjR7+A4YOfgIs3MHl1B+uf/nsgx5i/+z3svfQ3iBhg83N/gNmrf44Qa+x964/R7e9h8PDncfS534GrCoDIjObCG9K/O5dR3/sU1p/8HKrjZw6xkegpsyuYvv8OgAr73/m/EWdjwA1Q3/Mo1h94GsP7HsbuN/43uKOPYHjPaYTdi9IX169i8PDnUQ+mGL/1GpoL38Pkxnm4tdM49sV/AtdewmR3D+vP/R4IjPm572L/5W8gYogjn/sDTF79c0T2+Xke+TUc/cxvr1DFXUpLU0MOI+46uLVjWHvyS1h77JnepK/OPINjXxzCrZ9GdeREjwH98cdx/Ev/DDQ4jurYqT5zrp/B8d/6T8FuHfXxe9Sw9rNTd/UtdOMpRmfvw/iHf47pudfANMTm5/4x1h55CvO3vg44h7C7hdHjv4mNT/w6/ODWao5fPw6qh3DrxzC45xEMzjyJ+uQZkK9AYOx/928AtwZft9j55h+juXoR/thDOPH5f4TqyAbat4+i29pGrE9h8/m/j7WHPgZyBxmLI8OffASbz3wFg9P3fyDzkR/CbxxB6Byq0w9heOZxDM48CjdcAxGhu/ZjtHtjDB//DMYvfxXTd14Fo8bGc3+I9Uc/iebct6Qvdm5g9NhvYOPp34AbDjH+7l8Cbh2+mmPnm/8nmmuX4I8/LM+zsYb5T48gbO8g1qex+fnfw9pDT64ExV1M9Nf/9r+79uUvPn7qw27I3Ubzc9/Gzve+Jj9cjcHZT2LzmS+j2tgEoK7CZgKqRj+3QOoRR+x+6//A7PIlAACNjmHtyV/H+hPPwXmnh3SIzRxuuL5Upmov/ABbf/tV+eFqDO5/Ghuf/DLqI2KwzH0xBPnq5s/zsS9i/fFPLzxPk4TSiu5e+tYL79z4UJHF3UyDB5/DUbcODoT69EPwG0d7E5qIQMNf4AvoibDx3H+I+vI50OgYBqcfBA2GPcWJXAU/Wv6QVfc9g2O/ViF2jPrUQ/Cbxz64L3rPc1yfZ3BXPM+Kfj5ajdRNiPwQo4ee/eADf3F3hN84hbW7EOSRqzF88FM/61l37fOs6OcjB0gMQ/rDwveSDjuGF/YfRj/LOfwBn7d7zGHnLLb/Vm292Tm/iH45rN2rfrmz/XLYM97pfrmd85bVL7fT3ls+K6GSHQU4/Fke9E6dc6cY42bn3mz/zbbdiWf8ec5Z9cvh59zqOX6V++VW7bmNfvnQc0NWtKIV/XLQSlisaEUrui1aCYsVrWhFt0V3nbD4WTJgmRmhC2i7D06NDiGmdOimaRE5K2ehC5jOym39e/w8JOcx2qbFbN4dep3Fbcws7dTv1tZ5c/B8e54VrWhZtDTXaTtv8Obb1/H4E2cwrICXv/8Wjj74EI7QHFszxpMPn8B8MsE3Xngfv/PbH8PW1W28c2Efn33uIXgwAOplRjMDW1e38P+98A6O3n8fnn14HdcnjI89cgLzyRTf+Pa7+MpXnsJsb4zX37yEn5zbxj/4R8/h6tvn8eKPLuP5Lz2DQbOPN356DR0TuGtxzyMP4HNPncLVS1uYcIVHzx7FdG+Mf//Dy/id33oc7kAbGJfOX0dXjfDgmU3sbW3j+69v4zeffwA/eesS3jm/DV/XmOxN8Pkvfwr3H/E4985VHDl9AqeODnH5/cs4twV84Zl7cfniDfz4zUuY0Ai/98WH8dabl3Du4g7qQY297Ql+8+9/BqfXHPZ35Xl++u42fv8PP4sjA38wY3xFK7oD5P/LP/ryf/vIQyfX88uG7szf+ct7ePHl9/HoI/fg5e//BD94cxsn1hk/fOUCJtHjng2Hv/raj9HUA1x++zxuTDtc2+nwyL3r+Ntvv4X1E8exMaryNWPA91++hCEFbO9O8e5717HXOpw54vFXX/8R5tUA1969iHevNXj88TPYvraNKxe3MHdDTHfH2L6+h8YN8fxnH8MnPnYGNy5ew7iJ+MkbF/D2Ozcw90Mc8R3+8muvg9bWcPG967j37EkMvEttmO7u4dvfP4e2GmEYpvjLr7+B4dF1vPHq+zh+32k8/9wjePLhE3jrrUsIXYeXXnof75/fwrEzp7Bz4Qr++m/fwYlTG3jxxZ8CwzU8dvYIzr1/Az/9yTXc88C9eP65h/H4A8fwxltXEJoGP/zhOVzdbfHEE2dw48o2rlzdw+bJY9gYVnd07FZ/q7/3zu9MVVicWMcdpqHr8JNzW7hyaQv3PnI/NlxAtXEEpzeA7fEc569M8JlPncX21hhPP/s4HjxCePP9bVy4vIdnPvMYzpwYgYrrkXN4+KETqCuPhx+9D+vU4sbeHO9f3sdnPvUAtrcmeOqTj+K5T9yHjQHh2vYMz3z6MTz1yHEMRkN88pmH8MTDJzGsHQgAg3D8xBF88hMPotnbwc64weWtOT79ifuwtT3FM596GCc2Br1VvB4OcP3SNexO5ri2H/Dsx+/FjZ0ZPv+Fj+GR+4/CO6lz4ZzHmftP4tlnzuK9d69hvLuPplrDY/dvYG/G+M0vPoVHHziO6d4EGK3ji7/2OO47vQHvSFxWlcd9Z0/h2U89hCceOYW1Cri+M8czzz6C00f7UZ4rWtGdoPfOb0/pr//8v19KbkgMHd6/sIPT9x7D2rBKE3x/d4ztScDZe4/AFUlRzWyGy1tz3H/mKKpDkqUWabw3xtY44P57jwiT/R1od3sP45Zw5vQG3Adg/K3ru5izx72n1j/wWGbGlcvbGKyv4/iRwSofYkW/NNTPDTFbGS18t303+36b5zhf4eGHTuWIMT1n88gGNsuKdLpvMBzhofsPSalevKd+bhzZwMbmwvbFc3DIuQv3BYCjx4/gaLn9Fs944tTRg/e4yTlEhDNnThzehpv162L7Ftt9s3ve6vOwax7WpsV23ep+ZXt/3vlyWBt+Uf1i9KvaLz8LT9zknINvUf9Zv/+izyl/38rYf7OIs5/n3Ju142b77tQzflB77kS/HHb/j2K/3OzYX6V++bvMG9yFrtMVrWhFdyHx6r0hK1rRim6TVshiRSta0W3RSlisaEUrui1aCYsVrWhFt0UrYbGiFa3otmgpwsLynQ57VWK5rzxmcfuKfrnpsGG8nbH/RcyXxeuU59xsft3snJvd43bbe9i1fll4YikvGZrP1jAfz+HIS3FXcgARyBEckUQy6nYir99lH4jA8FLynhyICExeryHXARzgHFivwdB7wAFO90PO1+go+Uyy8hdQnfsjQxGZtSPA9ttmKwMI8lpGRJ3F0OMiODIImgXMcj7bMQgAGBzlOsw5w1Yuz2Dod21DyqzVbb1MW9a5S5wZCXLNHCfAAAjyHplik33HwY0HsoHBYKYi9OBm0oKKS0mbSI/Ol+TeMf3rce+jbIv0C6XfRIQHHshvebvzRIXrlNM2HIj2KqncV55zC4qhQtd0IHJwTpjcOfljEwyuEiYmL+8BIQKcB8OBnLxUVwSAV4Hi835ygJdPVoFDcGBnAsVeylsIFxMcTHrN23iQjzRxnsCkAoIDTHiQCg3mINudCpK07EWAAwj2PR56HblJSOfEKILFUvIttZ+Vw6xswGFvoi8Z0ARNFhomxGTCyhveKV1bWc6OPJRB+/eV4yOZMDukB9OFVbCU53JfxPSfR5954aqLz8zM4Cjix6UF7yZkfHorXrbjsHDsTc65eQTnraDO4r4PgkVEIJQIAsWfIQoq/qB5E8U2QwiKMCyji4gWtql0txvYU6eHL7eT/b8iACCbuDIxCawrY57QgiYgk59ZT+H0G8xwMGYVoUGcUQhzEEQRFxgymkBaYPQeIjg48ViW73QOpbaXxy98UsntDAIVU3jhHso8RP09dPBIQb3aT+UtHAAmQScH7kB5C4EOecbFm+gw9Z7hJnQ7vHyzYw85Zyn1LAgmJKjHmPYrbS32Cz8vsrENUTnAeQCSQCrvckAS8AHJmX9+kBj+6BKnfwuhkFZdUw8MSRjaABgRxAGIQQVLTMeaSmLb8/mHNECRHRkSIM7jW0DvRWYSBs1Txb6zMvjivVS2pGHOaIrS8FPavpiuIYIQpFpY77r5DfCpjZRnFbMugpx7N18/3+WwZ+x3E5fyZam0pOI3Zff4QmgonDKIyAwmBrEJEc7bGXAUEdmBKEM2W0XIVhhmUFohOc8DlcaUtUiU+hSDfkXFREl5BpYaum3JgjYLXDLuJAIi4OBEMOjiwGksVeWE2DaAzGCEwlKit/EMMAGRhNFuzUA2vuV3zkzYO5WLc7hg1pjlUmpzn5FtW2QUWxcQEhTtKjKT51+o5MaCNqIJ1oXzy+9ZNQMoFnP+Q8hYXoqwyPooICuSGX1EJyWQqLeOExRmhaQ2YIYkiG1EA4AKRBGIDnBRVxOXxi9PBha7BQNMYmSTgxk2bIAr8MqvqtgoGcMBHHpaHMOpoDBRryKWZDu7KOqErX/OAdFQBSkDi5KSxLSOvyOIaTJmJKEiRrbT4czU/672iGS4sNKDdNNzWI8juz673rWSugukOUtwYGY4UpvKwlJPUc7I9gjkBTHfVVHUQaFTNBIOxg/SFk4G5w9FWNz5m9oA2qofVa+NHOGZFAlEMHudKCoAKAJOVh4OMifhWIUDAHQQT4ZY2IlVZDu5KUUdeAeFF/qbDlulIn51vSKH9QcfMjW4fyyrwMhWxf71SmZJ6mN/PsgVsr0DGTMCACKzQP4FA2a6U09QHC5MoCqTiTeAM9pMx6c7FiydD+pfLwsXmcd5ybH7AKbZ2IVzZ5IxPeWpKCIodSqinaKyubTB0GH61R0nWl4imU2OGBnOZd2AVfVIE4tzZ2Spn0xmuvIr8qBbqQ7ZgGmdLYO3YNNYkdJhjL1o3GTjdF3hoqgVzCLNjdntdwyFcVP+Ynm+GS/NlRpjHvsCfVJCC1ys8LndBzwliwbOEtKn5+sZLXr9kFVSQQNmc2OOyAo0kipAho5sT2G7ILsemUtX1BJRVUjV7qz2ZVvJ4XiDeu1Y7jxekoFTHBZmHDJvh3Nm9Cw9JdYJ2ROStifLlMvGK7dwI2ABpZXDm3dQgnZlS23Dr7Iqwjq9M1qgxJBZoMhQcMHoJkzEhcos6l5mOiTjIqOvhiSmXDTulWpkeQ6QLU8LgsJUz9TG8nppcaHMlES5PUzCyz0OLZ45qUJ5bhz0vJTPZbcvkVdhS4H1xyHV6fVY03AOPOfSkcWyhIUJBEAX+6LzFpnV+sDwKukqBahFmQEEMDu1VwSdBDHBPRlwsz8EWwayrOYortWedM7TknoS6KNOvPBZ7ulD+ZLxSlclkI16i/3ZH1Pu34YoWTAOs1+a8Fj0MjjkqVOGkPXOKe6hJ/da1VsYCpRyK4Bfqjxi6CwWn0LlOIBewEkgMNs80/0HbtZHd3xI331YBs7lcAVxRggsa73j/B4Pts7kCInqs08hVtxJhZ6b9eFyJQIA8esTFdOIdcVTN56tdCmAqH+BD0Vqf3hEh87XhMbSElz2Nx8i48teKwQF0EeF3FcEF1fqw6j0CKQbLo69HHhA9VhcDgimNsh1+kimePbDpNcCUe857WT7rvsou5nlJE5nEh3yTAolSI39lP6Qf1tg8pLpYFDWIgpf/F4eU55T0uL4J2wXQfAg26RCpFQ9UAZo2blmcChuKAEs9h4PuW6EaptmLKOiIWXbDzxAadwUz8ivjhpyc2QBQHX1wxi67NCo7u4obu2kPii6M3XF7A/pErZ6RvGCLBieS0Y+PP6AkzpKYEGLt2DygyiouA5yE6LFeCxcqlzNZXXvK7kGhvPNKHnnzH4BRkK+AnhLtKbPQgDgJNaEzAa0oDLdTFvmhX0HePGQ34vX6z1DpuqAunTY3Dk4Rrf+feB8VldTASeV0RkRkUklJSu6AAz0UDIGIU8upxK23AZVH4zX2Z7WwKo1i2GCIbtRPZgKoxGz/v4VUUd6glX6li2YwA4pV0czNhbeDl4YDz1JoXm+VmkTIAu9h60Jxarci7Iy5syCKwVeAYAytytQEi+oH4eRnJuZ3esFnaqy2T6QVZv0SQuIrGxXiVAPLFLW35Q/i+uWDGjCxQRvaa/oqfKLtMjDPwu/3ozvOblO7+wqKnMopmAWB5d90fKBSGKPEIbXyeucmL4iJThmPiWmKK7U6ER4AEhAKUL2JTHpi7bI6gf2kIkqsQTCK5ZoFgEWya4a6R3tnw+PjGsXZg9zwYy9sKHiGAeQJZQZGTokpLgKJg3UYu1fQZjl0i0h+1A7lDIY58ukVXVBYKTzIeNaLMtFDIMeb5Ge6fkWUII0ZKEPLLaHkaIkVJW2/kiy4LDoUlAWdMDB/R8QrdkzjhYoypDKcitM0PJeX1jGWSQ3WJSnZ2dwoAiC1Q5xjsGWgKY+cIoGOSVZjCwmg6KqMV6EAUUJDKIIaPJZ0p9T7I3sF7UGecL0dM+PLuWV/5DnNIQBm/jCKCwRVGB2KhtYhX8EW8cmpADpY42QhOFwi9SlzBQl8/SFVLrkoUChF/ykY8blb6Lk3kxu1MVrL4ZqF/cUA3q2tZgQTdcRiXJAubX7L2o92avSv39fGNpxhvZ0O6uL+UMwWixHWJRWdBtYykE2OZDFjlMGZkKMYqyMFiZOGqehUXSAzj19e5egDJMGpj/rakakQkT0ZEoRiQBTGa2fV0CWN5wuoZPuBirUCgBJpSBofxXMkfqV03HGppkhLbg+CwAQgR0DkTS+ps+oZUyNnFO2jRQFmqpYMqdPbcywhDXEHOn6eaXPasTiCr/ItGU7DNWkc7VDVF7krHntrB7uUnW6Zwo+TMKkWBN9DAAcAziKF89VXlX6m6OSO0FLEhYAR2VQ58TSy+bPhz5zRIrRByACQyaGdZagC5G2ZMYJGyxzqzKrGqFSiFmiPq0hOunIjivUMB2iwx/gIygw0pNSf0vuh6yD08JZnFQNRR1srnEVtiTIMYUrpYmfQ78tB4hhaoGGa8NGJf9OaEEFVW7K4tgCqc4G8rEp4zOd2k9ZP6xnUqRl+m5evbLzsnBVoJWRTCEESxuH0/5jLKAiPa90wcYYIHa7Cqg8OAbEGFQoLTfieImJZPatSOTSDhV3apbKJVMn5tZJKCsPZAI6V0zv8hN9PTzHy2YB0oPdiiKSgmxqke376AmKWxMvCE5xbfcFRmlDKo5RxMEF+pAeXMxp0IVhYYEkINkKLNoxx1VoNqqiBlJ1NcH1JHBccp1nJtdW9hCELhIL+4hccU62C/RVhFLQaLxIEkwsvk02dJXTF0245mhSaUApOGxhBQDvxbYWomXxAuRd71Wfy6LlJJKVnRMV2usClAdv8eE5wUaJrwCILDHIpTh8qYxl+q9CxAIiU1J0OU2mfAsuhAjlSYO+IMkr60dLaBwKZAuV4iBl4WErYEIAvStSIetLhd30b6fzITOreMtS2pQwY2QQ+WwgVNZjVUHk3JywJcLEGNMX7Y3FvRfRgj12gQRQiLQkSFCcn5+nFBrJOGvnFHYZ1X96/UrIsUSIERwFETmtFhc5gGMHMODJia0IyPaXm4zSnaLl5IYkXaN4wEULfBkToSdJrIXFXbj+n5MKWExOS+4RknGTHOCsmpatOLI/FclJgUK9Rhagspj4H0niD/jU3A0du6wu5vFLSVC6ZB7oqZ6MKCc3p+7NOMOEinkOShtSeTHT/fvh3im5ivM5xRm9ZpWp8/K75HAUTN2foyaGLDair74sBvdx0V8ue1xsEdTPqAJCMm8dIgKYu3Q/56pCOOVQfDE8L9e1v7TiN955OCdMTsjl9UjzQ5zLQgEWqEWU6naCSM4lLxNLBYXiVpiWa98JEo6bEQeQ1RsuRjojjjQQPRmR1jrY6vXLTyUzcG97n0QNYI79GItkwCwYwJBceerCJRl9z8AiS9u2EkkcFNj5dw5oupk7VY6nolH94zgZEOXRoqoAnO9iC8tCW0u3pgBU6vUBc96S6qswYFHKNslcUrkAEMOTxgAVKo2ALCtBKCjJ+eVnSFfSoLxhIVbkACUL7cI5tyICkjBIzK2wn4rzjeUBSkDDoCelm6sawwxCAMNn/ZIjLKqTWQciatAFxUMbzQggeCBGgDK8lXtZJKfp2ybJf5kFhkUnMkr38EEMZcIxi5RSiyvYRlBGWjGzKMp9V1xRmURUhkKOJ6ie1ZJ0no5nH13YNmuNXreYjM74s5Bcdm2LGg5dwGS8j+2tPRw5ugHvPeazOQbDIWKMuHF9G9ZZn/IAACAASURBVEePbWI4HGBtfV37wBqu7V1QLsoPQRCiYggasNksc42IJAjMno9VaLHYgMDZLuK15mwPkt2ESj69FX8mwU0ffE61aAleMCLf8gY3+33geJQDdAhgLRrHbJOPtFCA6XVOuth8zKmYSNQ+dllg6D3EvFFEdWoplWI6adwARGAwAAp5aiUOMRMbFx35yy0w+ilYGW31J36xive2KYPYkpgAm10n5/mILGHVz02YxMMnTWkg7G02QZAFhNmu8uQ+PMCJitlmLY+hEYTqHTi2GK2t4Z7BEHs7+zh233EMBhXq4QD7+xNsbK7jxKkTmI7HIGexOIJYE/qhlIgOCT60iuYxTWwiAvk8/5ld1sxSf2nfgKXyPUqUYc8Xi2sc7MJDuvMDjzvs2APn8NK8If2bSih1H0aVgShWScs8JenE9DWqtVncpQkSJr01FqKRQBzBkQCvkza5XkkHnrVatVXTSrMfGbLaKunS5PzlI07CuFTNxECcBUiOhlRk19MdKK92yf1ZrPiwldwMxrYCZ++SeF31OsRSLo5Yx1SjeNOtLJBvsdJUnj+LaCG7Ixexkvxuug6+EmY0d3xd12jmDXZu7OLo8SPouhY7W3s4++AZABHeE2LsCm4izTrlJC/tX0ckNjPO/Sv/q4pj58U8t5yzuCELD8hp/dJ2C2rLEak9nrjDxPgQhEVPBTywjw7/XvybdJdiLuT0Ggu2WbjBgfstrKgKFamHIqwuqMWO28144RqH3uAuJFvXS8OhrlK68qeJDRa1DCxqH5c9Svp/AZ1tQArvAsghqTqswVHsIfE0MdsKUg6KQXMbQeoJAMAYKC8qpZEyPxMf8n3hqLSoMKpqIMPMEUeObuLalRuYjse4cW0H9z94X7rKcG1dhWQuYkMWM2J1RxVdyX4TH9o/xCC2GKMiIcxc9pzbZShFGmvoTFCL5S8dWuztDtOSUtQXXiaUVg7q/dm2JB5sn56Rq2K4hbkgA595XyszKcoo/dc6QzNMZLNGA1I3I+RzYe/BKGG7fOcCVt/9VBg002ofFz4NbdgfFtAHANjY2GjotmSDKsfQTqVDZCnl01w/w9euudi3ROjNE7tPfmVE6TWjm/7l+xTH6n29q3HvfafxJ3/yTdTDASrv4FwF72s450HOw/kKzlVwnkBOVBly+t3JO25c8eddBUcuv2BLVSfqPVN/AbV9KPabgR+H9MNyiJaTSCYLhw6qTbRbPGzPfoF+R2bLfEottTskyOpshSOT/EgrHFQ691WNqNI+T9WSUYowsgMacA4cvnvRRUYUhSBIO/PzZZtDFhy5cHKxz4QvgBQ1m4RqcR3rI7b76Jiq+mECnorvBabX++drlyu2fC2yiQsX1mLodv9x1djoqX8N8rKwIGLWtOJ5cOhdp+fC5IVrc9nufEy/HVwcWhzPZfup95ypS4v+7RuQl0fLq5RFpG5Sd0DS598OZVq4oQqjA+t4skj3V69FD31CyTfBUSlP4FAVSQZZJnpxzwJ+350O1XJtLgQFL/wuEQbn75ZnQT0EZnUztU9SKT0WtYXzuWwvF+Jcp1NkhhxLJbP0ECBSO7N3Rbf2GPYwAdEfhcMEBQDEEAHXwdlb7FJ/icfizL3HMRwNe9fm9Gwo7mOrGlDGkXAxN/rtyMvOZLyL9fWjsq3sB5h+1te1c70OQx7LtVkAS37JEIDy+WVfEhiWHp7PyVARmZENwyVERNnd2buufdHJ7LjQgaUhYigSVCFb1VuSIvGy90SMoqmGs/xOuSUAwyUU82EZP9Nq1VM19HuBFg6qVFkgiLHT3iImRXi5x/QmQLQ/C6QhwkbLGEbzgKgQiLbfgrmysGAtmwjEXuEyLgVMsa33zOnnwT4vPSScCj9DFi0A5HxWUc274hyOH99EXdUoCyKJjSSvNgezRhfaUgDQHL6ui06qF5LdqGkuH7huVgHz4sdYtoETWKKBk8jBacCV03eZepUAFqgFmGApBMyCYDDJy+ZetYlKUGeFmToDAI9kRY5FlqSiGHYMik4hsQdclNoLmhFkE0xUFlV71KCVNV2bQAGmy+d1ZBlCgxf+Lf+QmB9A4fHIpQspCQpDUCx1Tdn8/GbTMQShn7YNGVFAvSTE+r4Lino7Eza80Gw1GGasLR+FkGjmc2k7gBADiBxilL4era0tMCnyfFlAIQlBECSgqSfQKYWam8ocNCZCvEGFsTY9Q5E7RCo8UmgAegtTP12AAHLwvs7CqxxOq+mCLJD6aU4M8fXbhF8eLSk3RP4tU3/lUVXjjyJBUwKPDVJPQGRDj/yp240I5iolspfamBDS4U8h3g4IOeSbotS8IKt5EeXFyvbiZElWi5DEJBUMyWNiSEIlvxmiCoiaICsVxsBfZI8yAIq9bdnWIMxs01V6tHjBEjMs18aECKX4AGN+RROA9KseK5A4ovcmdZQ6ek4EI2LAa1xBKAW27Jd+5tyPC70UQgcOAcP1DcSO04yo6jodXXjJwRwRQyeo1Nv0VqbTA0MM8KoSSwRlnykdOSmNgGLlTwiY02Jl12aG1F1hLFzLpF/xRJynsHM5fyUjD1o4TU+IGsRltpEPAbwerMF5B4iZEQODSL0LBPRzPgJk0LmwDJc2jew9sU9KB+YXCbGpLU6rYEU5hk2QmMBI3/UlRVF/O68vVLbsVvkj2DkW3aVMoveXCLyi5nTSm+Q5gMLNSCXe+KARt1mR2SiZWtNk5OJY+4wqT82+ENOnHKbRqgkd4MBK3GuCNZULUahFgzhl9EJXefuCQm3TTV5RodksUn6JPaOphnYfwsbmUTTzCULXoHI12naKUdL1+/kYXTNDM28wGK2jCy2oazAYbaT2AIQYAxx5ifdzVVINhM2V0Z3T+Uro9b/ZRSjjRwZUVchCyyKK03UNkKZr2FxmkPdaUoVV1TWBY0JcO88xurbDZDzF9WvbOP/+FfzBP3364HjdQaoSNruDxCxGJadBN4LWbRaWIdpBJW6RlEzqXzYPR7omF8dBBINT1cHCcdnccpqZSgDByvsthM2yE8ObMyawEHKFnwy9TpDVpUQWZCZSl+6VEJFRER6cC7JkhNC3c5jl3yaiHVv8LSQz2VvdYHc1tKDHJsZKJyBd1aA3ki8/Nbp4hmIF1MMFOTj04x8ycpRrexVxel1ijYS0I/L9CJQFTuozYDjawHw6wQvf+h6++JVfh3NeV3MLkJMrDdwGqnoN+7u7WN9ch69qxMiYjSfY29nF/t4+3n37XVy9fBXra2t44OEH5bxBjc0jR1CPapw4eQrEjBBiSlHgJJh1vHvGVBEGs+kY16/dwP7OPj72zMd748nMiBwQo7xky1fqgq1qyTAFp2ou8tgyxm3TYufGNs6/dxkXLlzBu29fxtb2HqbzgMFogD/4p5/A0oiXaOCUzNC+nzgjBvssQsJTIFRmPEorhOzv2QTsqyOUm0090Km8wHiZY8jJ+gsu04qV7Q2Wk6yovTqe6RJmCNXGGIREgX4KOJvKz1m7elGnWSDwArMe6Fsy24Le1lQCW51Sm/qPnDvNkEpGKf0Yh7wq55qUilSsY4kgrsfiGj11CEVfSWeXRs6UWEVZ2MmaktsxWFsHOw9fD2Ghzl3bYDrex3i8j+uXryKEgNlkijffeh9n7z+F8f4+JuMxZtM55k1AF6LNJOxs7+PChSsAo/f+j6r2uL4zxxuv/AhPPvEgTt97D0braxgNhzhx6gRG6+tw3onAgmSNdl2LP/2//gw722MMhgO89tKPsHlkE+ubGyBHmOxNsLOzi/H+FPNZgzNnT+P48Q08+uQTWFsboR4O4LzH3s4etm5s48qla7h04SouXryG8aRBF3SBY0JUsXL4bLiztCTXKTRj1PUExUHXaRGAYkC0JxTU/WqCw7BeUkscslbr0ouETOUBSpaj4i9vKZkprSA2yRVlpPaYNyS9e9XSlwXVcLJYxwP36hmnqPyyMA24f1xqUrH6JgtPkZMQQ6NMKHYK5ogwH4PIITQTxHaGdrKDGDuZ9F0nXgnnwCGiGqzr7SM4Zq+IrbLp9YMxKASXsXGuhvMVqsEIVT1APRjBVzWcqzQAi7X8XBbfqUp47xPpk4Wj4SuHd958Hbvb29jb2cON61uYjidSGIZl1QaA7d05YpiCQ4B2B7x32N1rcPTIEOCIrlNxGhmukvyhwIymDWjbgOs39tDM3gReeRPmZXIErK+PMFwbYX1zAwBjsjfBdDrD/niGGBnzpsPu7hjMV/JCEmUuBZbPndffBTPwwt/+SGZq5dF1EW0XUgg5R1JEIjPaqt8TJFHC3ywO4A7ScrwhzsH7hXoUhUHQBIUs6D3RsCA4imAu0VeyoEjHOrVR2DY9loprlfYLPY/R/51aUFzbGD6vQ7rNKXro8XoWKlycARQLfA/c5KCl9IzJ7QcAZlC0kOMIjh04dojzfcRuim58FdzNwaFDDJ06LiQiNRpjM6TgsWKhlOHIjBi7VF8BfF34NkbEonITa6o0xyAMpp4VRFYjKAQRqYxzVobAVxiubWLjyEmMNo9iuHYEVaVQ3FWpQ6QLA6b7O5iM97B74zq2rl7G3u4eXnvtPVw7exQxMEKnyMlJGYMYIyqXkZ0jJ5qlCngXGYOBg/cEZg8PxrxpMRhWsOrdHk6Yk4Co710VQYX0guadvSl4dwJ3dUufUcYo6nxN9kcCoiU5soMkOmZEK3Z5QuSIZt5lDEraC1oU2YFgmdYipyXWg1KpyOXRUoSFIwfna61D45VvM/ORConEggtCRFbUAk04Y+KC2dUOwCpx2bmeYLHVT5i79HhQMmqa8JFhyEV1yqAtLmwPfYOnLflF1GiKfhRbRxkSyMq8iC1iaMGxAXdzIMzAYY7YNeDQArGRmotpdVfXZ1ItxDCWwte1JWCLMszh7gCBogqO9F9uj7Q0P03/XE6CIkbzopg7VFEHVFgUwqXjoCv4DLPxHravXkTydul8qAcDER7DEXw1wM61S9i+cQ0xMkIXESIjxIgQI8jLeDhiraTFkoruHEIIIJJ30HhPYOdkH7PYzLyH917tXRFNC1TepbEMmp9YeUIXAKe2lYioZVxJ2mD9RYTIeeYyuP9OrOgk6ZmQUJ/0q/zFJFFFgMMRHOuaQAznswvXQZCJV5uQ76mTyyET6XeUnAN8JV4FKpg2rc6Fb7mM95ffDpE4xcUbekjtTiNDB1CGXS85F81kYPoxU1YVksswt0kSHWOqO5AqgkPvyZAMWla7QWqX/qnBMLYzhNkOYjtF7OaI7QQUW8gLhGMWakBicEG+nJCKrTwJeXB5fOHJWNyum1gcIMI4Zlew/bFQX6xnk0bAvT97dABgZ0LKDJNAKqiqMLo8z5qYUrgBMHeYN3OM9/f0Devy3GJcNF8Uw0eHqvIY1jWCE7RjgtKQT8VOvBzewdeyDkZ1+TrP8L6Fr2RsYiRUdQ3vCW0rAsA5zWFyDsQRlfcIMWfdRnNrOKmJaYmyQC6qw8z5hVnFdjnMYjnkftGRXAOE6BWz6pwBS0kG7wB73wol4U/wS5cWtKSyenAAeakBcABFCEI4oGLoZ6lS5FgHabMs4DkZiAtVJjFPzHCw66Sc+nw6A8Bo24C2mSMyw/sKMQZ0oUuraWZkgd2D4Uib5rJQskpfvgLHCF8NxL/PEd1EBIS4MtWv77zKMpmA5KtcJcxlIZpsL4VMzKpNwgNIkLZg7rTSJwFi656OBSxiEoWA1DsWalSWuTY/7DO7RMUrJOLHab0H5uKQpFFpanoSEpzaqkg/3dcR5Yz2yqNiMSSuDSoMhxVikN8hiuFPBJ4TDwYTfOVQVWK/ctEEL8FXHtWwkvtFhpsHVJW42ieTBoOhFFXyiiy813IokRCivJ8XaVErYiQU1NnKTxC1xTuS5F1TREvVOwrz2bFQoSHyVsZehDilMqakcz7EmITUMmk5NgszXmoBm8T4pMC3EBSsx4vuHBGCeCHaeQsihy5EtG2HC+9dwPXr2zh2bBMgwmw2w3hnD9PJDMwR83mDbt6AiRHaBiEGdG0LwFYQD/IEVzl47+Frj0onmfcEX1X63aHyDt4RqjrHhqQygeQEGicDrkQIkvNw5OGdCBSnNUOdr0S4mGAg18uJs9UeatgiXelySUIoOnNqUMwoq9BMYEIn9orcJLnRX/VZdsg7UjTk25HYRsmpeqNh9xoBmqd2BGsthjLozgRB1NBmUbtMTeLEOFw8Nwqkk+xY2gfOeQxqwqD2iBUjBkIIwvQhIquhDNSV07GS9ZBVOJBzqCqpaekjy3gPavjIiLGGc4TYBdRVhXkTUdUeZjh1TGpj4NR/UVUuMBDIvD7yDF7rXZCXwbVurojA+ha9CkCI0sWeC5ezwkjvFSmpfSlEGSfnPsLVvb/3wo/w0ndfl4EOEVVdY3NzhK4Nau0ldF2H6VSCapiB8WQKDhFdJyt913UyeWKQyWGzjIDKCfN5ZxNLGFzMEKLfkid4hbbkHLxnqURESNZ4gtlTHJxev5k38KMBIghNwxgO6p7aYEhJ9OIOVV0hhgCKjKadYX1jA7PxGHAmgGpNV3bwVQ0iD1cZs6vOn5h4EfqnZVrvnmJgISDWSgFA7wE1LouASsVaTMNmDYoq7BIiuHTiajl7IpcYHklcKYPeRFUBoC8i0+tEgGWZ1qzgMimLs7xMej0npinTuH2lY+MdOHp0gTV+ISI4QlBkQAAqFWIRDuSkgI3BegKJsKgrEIC2jRiOKkwmIkRE6Gs8CAVNTCY4dmosZniWZ+xCBEXAJ2RlGI7VNmHCUGwQ3rskEZxXVQlA6MS967VGbSTAqbDaG8/BDGyuD7A/aRCKPJVl0VIiOK9vj/Gd770F73UyA+qQMGNV1tt9skEARBYWTvBquCrPY4qQoMBiZVVpH0X/QCAWFBAZkSQwzPmQ7CeIBHiv23WSOML+7hSDYYXL529gfXOEtg0YrQ9x9uwJDAYVZtMGTddhc2MNG+truLa1B+aIwUDUiroS5CGuSdGjcyi1MHIdxegW4bW+oj6AMnCMBs5lJU+Rgaq72sDFAtqHYoVO7yHVxKOEinylSCivlM4unMiURS6yeKn3LcVayGCJ7ab4iyHCk8YjUNC4NNL22bUK749IoJ5tJt1RUahzHuWiWkdoMVu5XwiM4bDGoK7hPRJjB62KVQ9UDQHDeYdKbRhV7cUmMqwxa2Q+VlWFGGXOGKpgZjjm5A5lMGrn0HVcqGGi+uzszuCcw/r6AHvjOSazFrNZwLEjQ4QoY7q1M8FwWKOuPC5d30eMwNpQhHvTinE4xIhWhaJzY4QADEbxjvPtIlXLuKFYmEUSBo4Yepfemi2b8wQJTHCO8zwnERoBss2bRm+Tmxychi57e0OWY4BlUnnnRPf0JIZW74qVymwCujIFmSRtA1y+sAXnHLouoOsmcN4hdAEXDOI7oBpUmDcd9idztF1EVTm0bUBVycQhR+jaDlXllbnFYi95BA5t14ACwQePqKugcw7kK3AUpGIeiaquRPXgHPJ9s2zMJDRte+EeBYCGc5xEMtxBkBccZXdnKg7jADIrCmX5AG2LIZMFZExqACXWaxYqibTJZSMyZ98M66VMJbOlILl1yeaA0zg/L33qHVyIGA4q1LWokyEwootwEagrUqSpagkBXvMz7I0RXj8ZjLp2iNFhPm9lDBxhOu+wszMFWAK4JrMOe/vz1L+zRuwJg8pjf9KAiVB5wryV9PfAEdv7YicLluO438rzQYy1TWhTHLAZSQ37dUGqAdBCXy+DlpNIxsC07XBtHNBGxtGh13KLAtOGnrA28Ki8QDkXKBnXnOZ8OGYxYEYZNNmnSMDcZWoLcN5lFJJsAwZn9RgnhjDvXRIgtXNw3mFne4z5LMB5XVWUGUJgzGYNqqpCPajBkdG2jBjn8HWVoLLc0xhS7C/Oe0lLdqw+fE4TFoiIGm4eyIG6Rg1oQNs2ULikJeAowf+D/azTi1WlKQ1wnJmaCkGS1J0Y0QZLNEP2kBTXTZ/6r8Ws2Eqf42VMSHAKorN22Hh482Jo6HyMVjIuqyGkSMMiVCNHhCB5RAyCc3KOIVV5FMJw4FEPPLyDCNxoxuwO3bzBfB4wm7fY3Zmhaztsb00wn3VYW6sxnbboAGzvzPGTN1u0HWPeBDRth9p7zNuIyayTSlkobBcQA2fl5HM8beFVqE1aTnWjCaTHG1JRIyrnWA6CCPCgKFntndAoIgAZNC6PCFV299056nRBmMm7U7AzE2u8rRoeBJpKUM1aTdgcehzbqFTam0oiAsGZW5wIYIJ3MqkqdXs5EyRmo4AMlHOUhIIZiJwGi3GMuHJ1FxubNe659zjGO7NsA9FJGAOjqlWAeamlGE3nT9moRVcmg60wI2lMAJUPbrYGjslQBgRFOJ2s6MzplQaxa8VA6gUBmL0g30630eI9kA2VWvOSIHEIKWbCuWSALM5Kq1rXtojaFiKnb8sqVI5oSEG+R9aVNESJRSBJJoRpO1SYShR5hqiITB/IKzpjlnENXcTO9hiOBDWMJ3M08xbeiyckdBHNvEFVV+iaOZomYDppMJmIgJhMOrz/3hY4BITAaAMjnBchRETg7al0EYD9eUDXdrLya7dMZq3GqABdEDSSvDEKh5ogNowQWVAtifDoGKk+kOGlqOpMF+V6cIJsVB6KQ4n6tpBIVOSRLBdeLAVZTJuI/UZ7XCcyk1WFYIG45NBGBrcMRsDxzRqVU7eR6oVEaqCCxU9J0Ev5m5zAPtHJZXJ778W45b0KDMiEChHTWYv5rMX+fovJtMV8JkxQ1+LLJr2Bcw71sMJwVCfvhI2VZRBmm6twga0sOvtFr0+rbBmpaT2VYToBiFoUhhmSFxAjyEU4fRM8tLK5VTjPlhtBIllVUbUFtlob0lBzJSFBfEbhtTAkEQPmbStCDySoinPTxcCIFCEaY0y4xjlCDJyYqW0CQifPFSKjabpkYwltSLaHBL2DCGUJpQ7Y3Z2i9jIekUUARYYYlYkwHNZwrsXuzkT7E2g7RtdFeCfoMCAjQGIxuLaBEToZu6rSTOKYvb8Wem092Wq0KjNrujtSbElEXjsadXdkw6csYub+rAdOA8PkOaqKQEwYVMCwEiGxNxOjvidBG2sDh+lyS1kAWJKwCMyYdyy2BZiBUju0YBhbCOcd49LOHOuDCqePivHHAapPi4PPub5Kkb+LnUJsBjKQzveRBByhaRvcuDHBeNLovQVG7O13qCuxcwhAFuu68+KSA4CqgpaGh6IWcWlaDhsRqaqkrtGFV/cxmd5/uM3BVDRDC6yYk5xcK3StFomlNMmSoaIwMKKQRSnQK5rbkjRVXI3MTnXmtkOMQeMEfHJfWlNdlSNjm7ZD23YKpQkcsvIjtp8OoQsKaBjzeYsYAuq6EiQQGdPxDOSA0WiAGCUNu+uEE+pBhVbf9VnXFZomKjOrF0QhfDMXNMYgNO0M3jkMh6IexSCdMxwQWie2jXlDiLoIRQY4ABUBrpISzQEASARgp/3lUpKjpP8P4DAPUheDibAx9NJnBIxqj0HlEcBo2oh5G7E96XBqc4BpG1F7gCNhNBB1XBAKJ6E7aQNmDWMyF3SxO2fMOhmAyhEmTZR4kSXT0uIs5iEzQ4JRrHpYqV5A9M69GWPSNBgNCKePDgrmEwXOmF8KsQhUqyrVlYnhq4wkfJVjFMbjGdbWB5jNWkwmopM6B1SekyEUlI1K5hol5xBBoGhWaUUQ5sXRGBKzW9jqbVo4K8el1T2pV0h4vHyrd3K/kRgXI0d4VJCX2HTwVMNii1PGvEUPF3EPZjsJXavVzQn1YIR6MMB8OkbXzGCOS2agC52MApO6qwHAwVfi9ubA6GKLCHH1QWE1QYyNXQRiF8EcJE4gRLiagC6irj2CqpZV5cCtvDDK+wrNvMNs1qT3eBARYggpmmPetIoyxcgXAqtQiZhOOxWIipCIMGvEIyVdLcZEQCC+c4QAvT4Bg6GkvHuSpK4QJDrzyJrHpAmoCOp2JeyMW8yaIIsFHEa1w7SNmHeCioiB9YFH5ICd/Q6BgdEAGNWErUmLoSe0kTEPwKQJIvB0woSocSOQOdepmhsjo3YSWt5GoA2M9WrpRoslCYs0oYrJXZhzFeyq/13j/SGCY2/W4eTRkaoPwhVkBh8HDc+VgQSA8aTFYECo6oEwDAG+lriGGDts78xw6coeQhDmrJxDXRkSIXgCvBPduaocnCfUtU+qhoVaOyfuNgBpQjrn0sAbAwEKdxOSkD9ifR7LeYnJtAeLEGWOCDEk1S2E1qQpAlpQkHAdZjF+St6GvlEtJYCFlM8BnXiu6tCN54hdK1GtCPBegpe8BnnFKLC76zo48imqktS46onghjXMRcosRkSL0mUw2k7qk4SuQ9N0ScXouoC2i5jsz9CFiEEt0ZghlDkvEW0rAiF0YiiNkKI0XdshBKinSEx+IUSB9yzxFU0HdCGg9hJMNxx6cZMyIYSA6TxgbSjj5SsP54C9/TmapsNoWGEyI3gPQU4eCJEwbwUhDwdSIvLIOmEyi2gCIzQRzgFtAJrtGRwB8y7nmTABNRHmIaILYqOweZ8ikIH0fl7SbOJoC4J5/FR9qpcPLJaXom6YOFVGYhUfCsNUjkCEBvSP0HQRl25M8PjZTYHF2q1dCCDyGAzFzRi6CF9pfUaSkmujtQGGo1o9JISLl8bY3W+T4VRcqaQ5ZYpwvNhBZHIK7AMR6oG9I0Lz0BARI1B5ESS+Uu+KE53UqVu2fGl74vpiJe9pI2p8ZLM1qCpi79aIGlMs54gubFmSIXQpG5SttGCyPRjaAAgRzXQq3o50n4iuV7lbXLxitNQ6W6rGSGi7qBhdG0COERRtBY2udRB02LYtWrVDSJM5qT9d28A7oAuEedMCTCkYKmrgkvfCVPVQYGeIEV3L6LSQEjlC14hVwTkPJmA4EBVF8kGk1mbbSruObAzQBcZwUCFMGnAETp1aT9GQdeUwHreqekAN54JiIJO6GAAAIABJREFU9tuAphObgWMP5wPG04gmkj6X9HPtgFYjLYnEiDprGSNPkLfe6cKh6nQy4IMxD/YdmqZQ2I2YENQ+FZlRdx9RZKEaNywUxyIOPWVmEZ0/qhqQz2sC0HSSA9DMOlzemsA7wrSJqD1hY1hhfa3C8SODhAY8AWtrAwyGPlXRaxtxkQkCIDV8qgvVi1HUeRVSKlx85SWfoPYg7+WVd07qdDp9m7utTHXtUXuvz2EqE5JNQL7npCToamIGgWyzSHnW2lfQStBIqoUDgQKDSAsKq+2BY4B3+g5NqG5H0JqSHULoEEKAxW5ENQAClAraCGN3iJxGCeVbvykZYWNCFV3HaLpO8iM6Rl1J+bqujWls53NRaeraJwQTPVBzRNuQRC56h7X1GvN5QNtGVJ5QD5wsBN5paHQEd8KEoh5KTMNwWGE2k0IxQFTDakToRPiGEBFjA0dAM5e4Bu8J166Pk9uW1OjURgDEGE+bpN5UDoielIkZTcuYdoJubMEzdGtRl4CoTI4IHQOhFbepecXaIJ4SsOXGMConyLaNQLCQ8eT1YLRB7t8t3cBpiWQHXgP3i6cMupDUERA09t2gexYU0jwxMHYx4vK1MfZmnYR6Q3ValvdW7k5bzGYNjm3WSceeThvMmwaj9RE4Mq5c3cOsCaomKI8mphZ3lDOmVi4uTAuwojfMEZ5klXdwatXUlbcosiOzTFUXRREOeZv4z/U7FYlvmoIuqpucLe5Dyzzk1JtySqeuSyliS4DGMqjhLMbE2F3bihEycsr8jJqlJFXQJftLakFmNcQEBUBwyrzi8dDiMup5yV4Mj64NYEhEZdTU9qp26ELQlHPxOjBHMUSr6jObdqo2MZoIVRcl+pYjZ3QSVLixqCqSFgB0+rZyiSyXdlkAX4yMNoqdomnFw1B7U5t0wSCgdoT1mjCZK1qoCDU5VB2j6TSgC+KdcKoKd4iaoWoGbjHsi+BkhCi2Cu8Irb0tIRpXIC0ojmwxBSrHaEI2xIopSVRYT7QUvi1puZqPvcjY7BcomIk06IrNG4C0yHaRsTXtwEE6i7Xh5su2Y3YnAWtDgqNO9xHIe1y/McbWTgMHc71ScrnaoNXOJZ3RAxpxqKuFCgPxOkhUJwxCioVKV3YGqcek8AsIrLZoxmjFcxlW0j2Hdfcp2gwJoj8bRGeYKiTeFkMcXdtqbIIIrcCQXJoQEVWtkFqQKkTU/mF5GkSiWllYs9SSUFuCMmnbypjFGNGGCA4xuaklS5NUkKjBkaPkAMWIEIQpmlknka7epRUYEOTUtJ20IbCoEyG7cavKoe1UnYHItmYutS7aDqlStyeJyWAwuk6M3ZEZ0yag7RhqMwazJHJ1gVF5wqAiVOqejGyh8RGDCpjNYw6iU/Vyw0sqQggMBHG/puAqQ2wkUcqVjhc4q9limKNk5yLIPJ51gjgIBE9ipzCto9VxWnphPV5aDU6D4IYskPzRTpAdPOcoTE3f19XBJp1GsnFmdEMepH7sEAKaVmwGbeywPqwx2Z9jZ1eS06LGXYh7NWEZgBy6CAy8GBwjREgY3nEMcCSEVBTCAT63yxk0J2EiB1JBJ1mXHhAbAVGuTQkZ9FS4lg0x2Wv0yJwkyYhphVvEnJF/W68ys2RitnNU9QDeeXRdh661/AYx+sVgsRFBPUpm0BRXoCOXStWBzUsSU3AQgVK90ghILo6W+ReDpMV4IJ3PnF2cobO07IjO7CoxppgJsEVrsrzCBABiFkIxSmj9vAnifYmMJkoMhYni2hMqRYnzFqqeCPQXe5Os9sNKJuUsRMwbQlWJHaquHWoPDECoNQEtBMaNcYcQCV1ktACGlczfLlr4tlZbceK1CFFNFT4vjWJ3ACovLlumiBhle63ekhhEwFjZCorZa+g1eHHZtLyXDEFStxxlqy9DoFqlxsAIswZLhzgH7byIEFyK6zeVfDRwGFmGoCKAoMVDhoMa9cBjMu/EYKWQjTmjCV9p+FQUnVggJ7JawGovEIc9yBOAXKjVsaoHBVMka7baIhBZyrsBAKungk3gmKBQZMEOEQKTswFTDY+FeiRR5CJAnKswHA7Fw9C2IDBC6GS2ViZAZ/DOo20F4nedJJxxjKgrh8idrI5JOxY93HtJoIKqXiKQBW0gQvpDg8hmsxYcI0IrrssY5BqtekHmjahXbSsCmVlzNpyqH/MogiYgqQzEusLqItJq3UxEMXB3QXKNoqp8jkQoMAjTToKeRjWpN0FWde8YHEW1i5ExbyMGkooK5yWSdDSQHJ/AIgDb1jJ2gaNrDhwFRTSpH9W649TLoYt+7QEXzcMn0yhoyKcjEVzy7huxY3gi1Op5qZzYPkzweS3eHLVPuuXHey8vN4QBdJC6AObpMDtBSQFABUnldSQ+am7EC8FqlIoRKXvVVjBPpPYMrVvgxKi1P2kRguiXyQsTGFy5VJik0oKtDupaJGGbECNcJI04lJXZVxbmy/mFLwpnQQFQ9QVM6W1nkSN8dKpwCZG+rYtsm3CBwHJncR6mxuhKrV4AJlKBIpGLzbwBHBA6ibIMsdP6HRWaphE1ogLarkuZmTaBuxDQ6XYJlhIm6kJQRChIzOIPQscILaOuPaq6wnw2RxcC5rNWs04hZ5HaG6AwW4vkho7h7IVgZqZh86awnlMiDEVNjhO89+pxMMQiCbiiXgzJYd6J14EBzJqICJkPlnsBiJdrVEtRm4EuEGKkZFlggua2kKA4R9DIYEJdO1SduInbyIiVoFFLZ5DoZOg85VxqD2IPKZmd7QSwqjGkiZGWLyJtigS0nfRbF4EmfESRRZKqiSuypFZ7JIoP1fGlsyeNrPZmbDwyJOzOOMFIuQij6cSF1kWGm7QIUUKi96dSB4M0+7Qqw8ZJArecekgiA4OqUveo2R60ZA8RXOXzahsYnWNQCDKBDDIpfGYpRgB41krMZogxe6GteIAlSxnTCBPoZ2HMtHgM6Qu1g4giBuoiggZRhcjgLqrRTaA/IHEQlrtBRNrOkAoMRZbZSFp0KAYZFeeA4VAyROu6gtM4FDBjPuswGHjUvoavSBO9gNFIQsJn00bURU+YTgHvWQ2fUVP4pV2hM0EhkDwmQUAARbRMSQ0yVUMMs0ip4d5ZfUyHOYvBsQ2i0viUeSdjz/r+ksqLnSOqChOI0QVh2C4K8vVqsGw6Ru21rigz6ooxdA51I9HJFYng6KKiBkUQWl89eTBsmXPICWQmO0mhVBeRksZmnfBLDtKSdi2bllJWz5FWj3ACQeU9mKpSEGOghUlT/QKtv+AVKnIkDCpxCUYGNofSjZWHpig7dFFNigwJngmMEFr1dqhFPRA6jqiduLLIkaogXuC0d5jPO0EvXiYzWJJ3AJbYA3WhevLgIK5C56QcG3tLepIclZBWWmF+YW4N1nJaFZsBK7ibXZmchIW93zNNDTZ7B6PyYt8Qw2OHGIJ6OKKGOYuAaUNA23ZikIwQoyQMEnOaAs1cgqiGgyrFjkhJ+oi5Vipr2jYdV1UVQA7TSasM51B7h8m0RegiRqMa62s1GISmEftIVRP296eIqt6EENF2nErkRV1lHUn/qYlBhDuLITKq9HTE6XtkKFcKJHGO1L1q9hxIurgDnGMd+/+/vavpkeQ4ri8yq6q7Z2a5FD9ErWla0kGCdDAE6GIbhg8++ua/4l9i+P8YPlqA4Q/oZNiCrS+KS3K5MzvLme6uqswIH15EVs/6MrChpihUHJbcnenu6qrMyIgXL15wE6sDoS3YMYoaF3da2cFbM6YWQ4r+D3HAGhiypzzKCGNfHraTL3oYxO+KOdvGSDE3P0izMEpVxOEaPJeghWMJU37L+/ahybl6QxzFVUCgUAluI6siM+n/qI4UR36cwdCSvRoM+afiDx9AUUGfzTtO0UhUVDiCnxpcAqQBL12AYswJkQCVIMdUjwJigTGVyTk76GqoVhFK46JAVmnNTtlnesYjjHZq0sM7AqQGCArH/6UllCY4x8ev5rwJz08h2pq7TqnyVg05Z8zTyBDeSVRVtVURmD4pqvkJXqlULYgyo7+XkezU9fzem03vuqRLTq5WUTUhJ0U/UCjmEh3GqaMKmhnKVHDYTyhzxd1csb+fmFrFRYM4kJhBNaHvM0oBZguSGH+t64A+J8zVmKwKQNZ4qH3zflUNwZ8FOGwAsG+qoQO2fYf9VDB0pE0vr+NrGiHKnOOgAW972uxp6lQUo4Pf1R11VDc6eDUtAbsMTEjQxKazgqXSV5WpRPbqTaTPaoLizM1wFFyVTNerR5pLenZeOxPdeznBFsn+5dStYPSRJZqneLJcDAJ4DhqoNzx3zKDXnhVAz1NGkHgaqTUuv0GRffhQ5IFQMu3MsZFOWLVISF7eY0lsIUMVht3eEajFkBKZhcPQQ3KUMs0xg+rVFe/l0NT6LJit8LoixzcDSvGN63hOSOkzOonr8BPXc3SkIH3KwptQhdagejN5DiIVHapXPir5K1B3Mg4SmLGj9mJHin1y7If3JaHvB4h0AHwoTmXKNhdiHl0veO+DtzGNI0pRqk9texLGvA0dZhgGMl+7PmOeFJ+/uMP19REiwDAkZ5gC80Qa97vv7FBrxRcv71H2Mys6/qzjv8nXj5qrkoEcCeIBlYxQBxhVCYZXByCji5TlaZIBQ71bY00iulCXaIXPi2SqrsqDTuMueSOiCEbfCgJBgaFP8KFDgbzxT7+89llmC64V7oFr+fcUswCidMq8PprGgvHUp9NW4EY8hBow10pAyLn0OSVqCbSyEh86AGSpMEl0BGYoAkAShmwsU2VuNBGvWytZgmThOV9BDRWhWuUXH6cVSF0eBmIXOheMDlUkEQxDRkoOciYBOp78GqmOO8EmyOMAaS3sTgTMm+IYcjA/dwDQgo/ilRYDajJ0XvuPeRbqaUjrfTFxKrcvMuXPQu+Rzo2RS/TmQA3TNON4pMBxFGvgvSEUKOcUrQIyKrVU3N/NqOp8Di97lqoYxxHVp23VYs1hROoVuE1OgmGT8fTJFttNxu3rA2wHXL21xbMPLjF0Cb/8VcYvfnkLgJ2ZgHmkwRRGhffV5ITbEM/Qv0eoVGnL/+Fangspr/VlILAFdqO6JEdj58KAYoJZDLsBuNgk3B0VXTYMHUvZfYpSMdPfcCh8VtLSjLZX3AmFOzDfC/EQKoDTibTnsvNMUY8ky95Awb1hbCZ4TWfgudjQ8RQ4zESDBQF6eWuyMmTrEnBQ87ySFPJJ+e8EsHhaTkVRIBj6hN5BrWoMKyn4q42uSxwgoxSCa0mFgr9qQEem5jhOSEnQe+mw6zoA5kQjRTdkFAfOkotwNA1NIeEnhh5PY/GoSbzsyEnf3AhMISQwDcCl9ZzGHdftK5ipU4vF2VXr97YqXDVq9jKld416VFEU6DrFNDGiC8ca1QamMqV1n3Y9yxpUO3cHKKxW1aKYiwOsha8X4TNJYJhPp8aUocyMjA6j4ub26NUtHjDXNwe8/OIOlxcDaqm43HX41geX+OTzPUrh8T9OFRnAcebnFjV07nSnahjSsn7MgLHC7ys8Gg0shPgIGZXLQcS0189/d+JxXzn6WXCcWUUyX/NdAoaeaTbbbS14WDw0xVXBnTFbjWmPCZype0K9kjiwaHGt57TuHJTRBKNeQKQggIfT6uzHwGyYAOTEMHDwwStzRWD+DLujfcJCsxMAhASe5ENelGCRKnCsBQBxD7OKkskbGPrU+AshB8frIxjF/gJAE5DVOFQnSGKVqNt4LL5BCmAZRSpy9jbn3YAuM54thUxJiDNOZOEYlOqt2gneebkIrbBRTFCKj8QVLrrMeJvXGsLGXukoxdWodYk44FgNtT2ZqpSZ5VEPPAADNpcb7LY9NqEvUc3BSaZ+Viv2e4KVUKDMBdNcm9hxzuLRR4IUBapfR6OZ+7PyYTlxP5miVCQ/9YvSuVWtOAK4HyvkevLKmOHmbo+5UKfiatfj8t0dfvD9b0EBfPb8Bh8/v8U4KY5Txet9QbBmzVipWMh+Cz4RTjhO+bYhHVj0bBB+O5ffQ9x/RhkGRipjAQZ/rmrg/TOm26QI0HkWBbhC4/Otpc2nFqnKG27kPGZnqoZkxxn4Sb6JQWBS/ef00gsVVo2oMnG6ODkdBPWHy3ySbr4mzmSARVWFC3FSbixxlpwJUItAMsuUQy/ttIvRAeLgZgKxDHEgyjzXnY5zk3sDqNOgpaIIw1itwGbbYRonDFcbACw5AobjsbhgDpx+bY0gFABYKEdXX61UBPPr8tOJ+bXXUT3FqFUxTZUsTg/77WSVGwAoHU+dFepNVrEhuswZKpvtgKdPLzD0GcdxxuFQcHNzT76EsuW7zIpS2JRVVGGzpyhJWsoV6uGq8FKstaoE6eNRKjbgpB8mJ0EpXso0cTDUoFZwnFj+vtgRH7nbj9gfCoa7Dnf7j/H+Ozt846rHj//4Gf77Fy9xf6zYH6maDcMDRxQsYvbCnHBgGL4hC0vxduIowqmas4EBvg+n28XPGaXNCpRoXDzBNwLrqF75SoI2VkCdQWwtbRd3D/Ap6nx/NS/Hn9HO1nVa/FTZ5KU0lLJh4wrMxUhYyUlaDupShM2FmyuXquf+aoAQHXX+gU+BMmeF+ofHaZGjdJvpDIoCSAapXh5VQ4mmAQhqVtemJJegVsNmO6DviOIzTFbf5NJep9A2XGieZgzbHuM4oZaKeTZsdz2cjtAcBlXBM0uu6toYid+5widQKTB0CbUGdV4wz6ziqxpKqdBCrKA60AlY4zQY6MiCa1FjyrhRfcok4cv7Ea+/POCz56+9imOAa02XufI9DZCcMI7HBsrCnVWtCaXOyGA3rlnzfv44rClqBWnrtDdGHZtKSZCUzVTF6enR+KaqmF5zjsYwJHzw3gWuX0948WrEFzcjvv+dt5GHHj/84R/g+fNX+OTzO5bSHZ8IqUa1hc8BLCkXrybSD4rQwIgTiMVhF56BGzxGUgSmYQCsArMAWoCQeOwl3tU/09AYy2qnP+OfMWryTYxCGm/kfHYWZ6G21IxDvJcLAujNWuNYCJhGDteBNWgIw7RwHCxuhr9d3q+XKKX5lwvP79EBD0YqhVfjMRNDedQpzdUjky5Tv4IkroTNkPH2O0+w2VAsR1JGzsCLz28dqDIkVeITQodGIEvYEm3BaATmaUbyJio2ePE7TKVgu+2RfKgPhICgmaJYMEeJDocgDKsAnooZ2abEI7wyokAMU+bNiHTFEGK9AMjctNIqArNDzrkTaJ1J5DJQMcwMOlbUKoDUhr9Q0NdQZlLca/RgVKUgLaxVMeK5KR5yJQRx6j9saovQnGkD+2/MBNNBcf+bO2x6wZNdh4/+8C381y9f4ecf3+KdpxvUMiMhZAN8IyrXENML5+FEKubpbqytJMt6SiBwakKQsimm+T1r99IWXCPWtRgwGjD7NZgwLZEHKQ5TFEUweJeqSIY1JxbXeW47W2QRC8FkoXrXCkyAq1NFk5I9uA2RlsQJFo+SHYZ8EH3Qoz0cNzNc7XpcbDq8fH0EEO/veXOO2RF0Xpve266d3/HONy6x3Qy4uOiRwLB9vz/icDjg/l7x9K0LfPObl/jyfo+Pvv1NvPj0FYZNh2kumCYuTi2KPiWKwCb18ijBzqp0AGaG8VAQrfkiQPEemFIqhV5cw5J8D3EJeip4sW8DmF30JnCDMheCigBUa6NQ4wSTEXDj5xCTBU/CFvGAjlRHo6htTPNy7cxoTosqklbiDga0tE0dtCzOAYmxCPF5UYKMdnhTRngGcyfHX4wycrSGi0cEIWhcDZiPiuNk6IZ7cECP4vmLPYaO6dVcFT3Iy5mKYHRNjOA9KNiKkIX3M0dZBKfXmpBgC7YgkcJYq6pEVHEatdBN8i8L0QqYPLuOmaeRhmd3KNFpGpGGeJgssvzrOe3M4lyeIqS44dzgBQQQATRWXZag8UaOxwWexFAh8RyRAbz7pEMpFa+PC6lrt+lwuc14ecu7q+bsP1Vkc71OsGw6zXBAM+HqssdHH30Dr2/vMU0zri43fjpWXF/PrNuboNaCeaoYjxN2lxuIKS4ur/Dyi9eotWA8zkip83khAQSqj1Ck0yiz4x2xiYQsys22w3SkAMw0ce5Fra51kAwpZdeCYHSRu4RpLJAkGLrsIjS1kbQIknLJJ6GjCTzBzO+5b9KU/d8qgddQG0+aYB1R+qrqLNV4qjEzVuhEBFClw1NoE9dtdHZED0Q07PHv5hs3IrAgJy3DDa1tbDtZT2wpp0P91WcHvPf2Bj/6wbv42S+ucZwVfU643Bo2PYlyN/dUvYrDpjH1PbpR7+mRGHbl6487NTa+OHa04B5o1yvtvntm0d4iSqCtFGrA7D+Lfp+IoBj9UOtj9qhN4ZHM72tkET5Q/a5N6sIhQiQYsrSrR74a1OdTJ2oeUYh7cTqUhPtDcfLN8oG3dyO+vOPpB0ekBfDNyltd1bzExs/vjL0SX3z2CtevRpgIPv38SxcaYRgMFbwqB4yjq05B8GreY+gzLi4rcpdw+LIgNDu7XGCJXZilAio+oKZ4pWGseO/9KxwOE4ahx3GacLgnhjEeCzUl2KVGJp+/b0nc4CkBw6Znrl0VmqgZOs9MDzgmj04CAqScEUpetVRsdx20eLUG8FJmJPLWNEjJm9B2ykEMMWUMWBrHqhKLKDOrQAEs0gFFeMh1QGcVw4VOOjZFGikrNh3gpU5Im8oWbxdLxDzK+vzmiO+OM7770dv4+NM73N9PKGq4va+43AAwaazf4wzMHrHEqZ8TKyax9lqbuB9esZbjMyHL36NTtuEe7kwcy+Q6tuX/Y2UHOhol23SycwSLlENQfxb1rHOZIFq0fqsfw+dvLXwEFrZcwPQSORzgbEM/6fw9omvU4GpDyoXcZS4iLdQCYHuxIkiyanQCAlKHcwK0FBTKTLe2ZgEIekjG8xf7ljNW9dKv62rOkpHNcDjMEAA313v0Q8Y0FcxTQe4ztrsNbm/3GKeKoeOUs1BvgnfNxiR2hQ/G6TJSFtRi2N8fAADTyPRCzRvguuRpibWoq9vkBjyaAZPfzIuLAZCM/X5sKYzFvU5osz1DP1I87cgDq0hwkeIklPxXp48np4B3WbwRbJHhhwO1ZNtqC8mLJ/GhJsb0z7mQ5pCwifMYrPmTaBZkFk8nQb3PACh94wZbVZyhWhQ//Y9r/PmP3sf3/ugJrq52+Md//Zjl2VIw9ExTx6ngdm+wSTA5AF8dVM3ePwQs7eVNSxSneAtLyrHf45BQjbm9aM5ySWjobOkzrW18AXzqvKffiGcTEQrfUDxd+b2shvDp84v1mSCdwJuEzDsHjchxl0B+rd/4OfLAZBgSb3CXgQuf05ASH3CGl+0ESJ0Tg/j2KGrIwnDYkjizjw5sruHNgcOoGOeRzqHLTod2kLVjatQZuzFr5Wvmqhin6orPPryohDIUm9dYLeHPxAfodr2L0nY+4OY4IXcZ202HV9d7DuWtrnJlgPRAHbUNRZ5LsFLqSdrBFOzqrQ0uLjdskktbjBMjFPFBS8NAmvr+fsQ4luZAmCv4zFMBxnH29vzkorbU1iQ2EeAsN2psBjMSsmCMEIvrZ8RGIe/DWoNVWHVAEwIk4++pivdvRLRDR9ZATzCaSScblAeT4O5Y8S//fo2/+ouP0A8dtkPGJ18ckcTYaySGJxeZTXbVsOkT5kICl5pg9JJ74BC+VNHkFd07ZPHxBxB0bU3z4IPfUvW0YamgOI/ixFHwdy3iFeqyYAFPYx+1ERH/3y35f7AOCK/3Wzb3sKFH4GA/fOkASJ4PL8Np2+xHoffedD61DILjTJl3nvz+u2o4zpRHa4CThI6jtHp2VebmSQUJCUVZ6hyLS62LYNLi1QxeelHiBVMFYAQvm8qUkSmJ0aB6xLAd0OWOszoMGMeKlICxFHTkSmNTO7aAC5AmDk/WWXF/XzHNilJmPykdXZ/9JG4VDsrSZUsoE1meKWUMW6Yk41gwdBmHwxHDMGCzGVz9nAN/j4eJJUtd+BxAwuFucs0Q3ufOX2Nm6PvBW/uJrfD0900OoJTqcnZoU7faiEMQUwhCXTxfpiPKHh+PmGbz9MVXB0lTQVYLZwG2bANN+zLatuk0BJ/ejPj7n/wGH77T4+b1hP3M6GtbFbteMM2cVpa9f+bpzmeAzHzqs7qAjUSKslQpBKR/iy34QzEeQAp4aTvSE0YTXrBqER48sggyoIpQi9TitZ6SOB7SUh0s0c05rTvHB5p/sy6zlTzUsbSFksQUkrieYeS6CKfCTXw/q+MU8FPdl7gQ+Nw4bjG5iApbmKUBnCHZV5Q07amBdSA/AR7RJEBMoT5FHKYYkFCchAUwVeo7Redszaqkdk+T4BIV1JvIOB4mLxvymicp7FGphn6iGlPXUdU6p4T9/UyClzNTDayikGjGe6V1mWvS5Y7y9N4QVYu1lEQg2F1uMQwZ08TZnUkE+/sJ+/3MVAa8V9NUkTtSpYHsA43Jy0ACutwhZ7h4ToCV0VPhHA8jhpSM+iKqFVXFNxTrw1qxVEt8w1SX0we40SPNiKY5AuFOivMoJiDO6muL/TIe3sOaavbPP9vjk5fcqNs+4dm7W3z28oDru4qnlz36juXQTZ9wOFD0JliYQ79wKPwqmOZYkKLiucb3YXThAmIOyxJrWpgVaLvcxE6chjRAk46U30WXX0HrRsCC45zN7IzVkGoEJtXQhEUCn6Kq0Ekd2ewNMIcLaDZmKCnAN3cyVdjKPit7ACJ0ZTZsyI60Fy+Vdska34Nt8ewXmYs3bKkhRtYRI0kt9y6VYWwKclktUAOGPmOqigzB4Ti36CiljDrNrXSMxJb2WhVz8hb2ys+7vBjw1pMtbsoe4nwRrUr9T5epyyk1hqRFWO9lvqHvsNn07AAdBnQdJfbvvzw6rsBUqRR1Ehlw2FeMU0HySKDrks8YYbm0c8EfVcU4ljY6oFZ4lGOY5kr8B+KS+4uzJ11/YS1y3xF7sHju7kxXlXIRAAADpUlEQVQyxMl7Dpi2DjZwNUg0zUVqEiestU0dDWW+j2EADrPhyTbjw/e2+LMfP8M//ORjvLidIJL4s13Gs/c3+Pkne2yzoo6GTW+43HR4feBW750EeJispa3x+Vnimhf+BgBGszBUv9eB66iYVzTIyBV/mgoyPeM9w+HH9witD/H3Predh5SFCKdZaw9JEvVcPqpS4Svj5GDvDctY1evZHGvn/z3x7NRSsSacm+AgaPJ5lWnpUSke6onBOwkVs7hIj/iDsHBeXs+35GKpDNFnAHBxFREBSpRmBXNhVYIUcj7UuVQuMtfPSCoernv1pxru7ibstgM2Q0/OxlGhlQxOqn1lhvN+Ck8TmurVMCR0HZu7dhcDxuOEY6EcnnoqVGppJ3it3OQxaKnrJGQ/AWG0tdt2KLVinmyJjuDS9k4nnwrp5TmjdbdOTgqLDTVXbVKFJM06WeukbAoEPsUXhTOJ8ztSllOeQjB8/Sk01m8spFCgUgPuR8XLuxm//vUrfPfDJ7i+u0E1wXeeXWI3CHIyvLXLOEzsHD3OFVOpbCUHnW5gKgIeTJ2wn4NRa0Q6guyLWWALSBo4hyw9ICRccX0kRBrFn5zKErzpFkQaxe6sdpZqyF/+6bfxvT/6a/9b4AB+1DRI59TC1/ricU8cD6rdeCyhWYBAEr/kDyneQzyUjBO1Vd1k+cR4n9MIL963aX7K8vnxWXLyuuTF8qb6hTg9H/7+6Ye2KdxgSXPhHrxxgba8zuz0mn3BJQ4YrkrQMyVxNW+CqQuj0/Uf/OYlWd7j4ft5sx+wOJI49T31OrU45eP+8QQ8CaFPvtvSKGXLSrCH73X6tU9/FhW1B79rD19n7X4Tr4qKxtU2Yegz/uSOk9NiBEBKVLaaa8w68ahX/OBqJKuHnxvr0t74/IfX+qYtD/Ph94x//987Aic/EaBNqTufnUkp69kHV3j2wdU5Pmq11R5lH37VF/A1tK+iArPaaqt9DW11FqutttqjbHUWq6222qNsdRarrbbao+wsGpyrrbba191IOMN5SzCrrbba19HWNGS11VZ7lK3OYrXVVnuUrc5itdVWe5StzmK11VZ7lKUV3FxttdUeY2cZMrTaaqt9/W1NQ1ZbbbVH2eosVltttUfZyuBcbbXVHmVrZLHaaqs9ytZqyGqrrfYoW6shq6222qMslbnuv+qLWG211X63bZ5s3/3zT3/2tznL33Rdd/FVX9Bqq632u2el6OGf/u0//+5/AER836hfEVzRAAAAAElFTkSuQmCC"}]}
