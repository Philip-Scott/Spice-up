{"current-slide":0, "slides": [{"background-color":"linear-gradient(to bottom, #51a7fe 0%, #022253 100%)", "background-pattern":"/usr/share/spice-up/assets/patterns/subtle-grey.png" , "items": [ {"x": -220,"y": 952,"w": 1136,"h": 456,"type":"text","text": "The Title","font": "raleway","color": "#fff","font-size": 50, "font-style":"regular", "justification": 0 }, {"x": -211,"y": 1211,"w": 951,"h": 297,"type":"text","text": "By: Felipe Escoto","font": "open sans","color": "#51a7fe","font-size": 21, "font-style":"light", "justification": 0 }]},{"background-color":"linear-gradient(to bottom, #164f86 0%, #773E9C 100%)", "background-pattern":"/usr/share/spice-up/assets/patterns/black-linen.png" , "items": [ {"x": -20,"y": 525,"w": 1527,"h": 294,"type":"text","text": "AMAZING HIPSTER","font": "raleway","color": "#fff","font-size": 28, "font-style":"regular", "justification": 1 }, {"x": 390,"y": 706,"w": 715,"h": 297,"type":"text","text": "Subtitle ","font": "open sans","color": "#51a7fe","font-size": 21, "font-style":"light italic", "justification": 1 }]},{"background-color":"linear-gradient(to bottom, #ffffff 0%, #ffffff 100%)", "background-pattern":"" , "items": [ {"x": -193,"y": 53,"w": 859,"h": 307,"type":"text","text": "Small Title","font": "raleway","color": "#861002","font-size": 28, "font-style":"regular", "justification": 0 }, {"x": -199,"y": 250,"w": 1924,"h": 738,"type":"text","text": "Lorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim veniam, quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo consequat","font": "open sans","color": "#666666","font-size": 16, "font-style":"light", "justification": 0 }, {"x": 1447,"y": -411,"w": 176,"h": 585,
            "type": "color",
            "background_color": "linear-gradient(to bottom, #ef5b5b 0%, #861002 100%)"
         }]}]}