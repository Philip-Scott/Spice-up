{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"rgb(170,42,77)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/inspiration-geometry.png" , "items": [ {"x": -613,"y": 599,"w": 1830,"h": 687,"type":"text","text": "","text-data": "{title}","font": "open sans","color": "#ffffff","font-size": 37, "font-style":"semibold", "justification": 1 }, {"x": -612,"y": 1171,"w": 1828,"h": 212,"type":"text","text": "","text-data": "{subtitle}=","font": "raleway","color": "rgba(255,255,255,0.59507)","font-size": 21, "font-style":"regular", "justification": 1 }, {"x": 1247,"y": 488,"w": 992,"h": 1107, "type": "color", "background_color": "rgb(182,59,104)", "border-radius": 0 }, {"x": -709,"y": -607,"w": 1958,"h": 1098, "type": "color", "background_color": "rgb(245,57,109)", "border-radius": 0 }, {"x": 1248,"y": -67,"w": 1011,"h": 557, "type": "color", "background_color": "rgb(252,186,86)", "border-radius": 0 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAZ40lEQVR4nO3deZgc9X3n8fevqu9reqbnPjQzkkASAgtxColDCJCNCeCDw5js4+SxTXjA9rMsD142JnGWxLve9TprP7FDNvbGT7yxE8c2EBuS2FwCyYA4BOKQBEJC54zm7jl6po+p+u0fNTqGGUmlYfpQ9/f1PHoeabpU9auunk//6le/Q6Uu+bJGiDJgnJHB+/vJYhejbBnFLoAQ4vQgYSGEcEXCQgjhioSFEMIVCQshhCsSFkIIVyQshBCuSFgIIVyRsBBCuCJhIYRwRcJCCOGKhIUQwhUJCyGEKxIWQghXJCyEEK5IWAghXJGwEEK4ImEhhHBFwkII4YqEhRDCFQkLIYQrEhZCCFckLIQQrkhYCCFckbAQQrgiYSGEcEXCQgjhioSFEMIVCQshhCsSFkIIVyQshBCuSFgIIVyRsBBCuCJhIYRwRcJCCOGKhIUQwhUJCyGEKxIWQghXJCyEEK5IWAghXJGwEEK4ImEhhHBFwkII4YqEhRDCFQkLIYQrEhZCCFckLIQQrhgAWuuTbnh4G631tL9/8PVT3d+Jti/GMed6/GIc82TvWyGPOW1/FPvannTzI9toPf3vc9lHPo55vP0V45iHeR4ae4d2y3/yo54iozqKTmfRExnwejDr4tiDo+h0Zt6PJQDDmP6JKCAVCqB8XuzkKBgGZn0cO5VGj44XtBzm1gDB92sKesxK4rE1zPfHS6NRhsK2bQj4MBMxJvuGIZub5yMJvB6MRAwApRQ6k8UeGp3/i3oihkLbNtpjYtRXYw2PoVPpAhbAobVG26rgx60UnvzsVoFSKL8PIxrE6hmCSSs/h6pkSmHWx7H6kuhsDlAY8QgqHkUPjRauHIYC08BsrMHqG4ZMtnDHFgWTlwZOBWAYGOEAVveABEWeqJAfO5WG7CQKhQJ0cgy0LmjFAsN0rnXPoARFGctTzQKnOjwyXpR76IphGGDZM36sk2MUtDJuWc6XwixlEeUjb2FhD49NfdeJfNHjaScwisweTcm1rgB5Cwv58ACGQkVDzm3BSB6eDFh2SXyby7WuDMX/WppPpgEBX2Hv10/E1ii/ryR+ocuOAhX0oyWnCiZvNYtC04ARDmLGI9iZHHbPYLGLBIDdnwS7ZOKrfPh9mPXVGLaNtb+32KWpCGUTFgrANJxn7aXUIi9BkRfKY6ItC53NoUFuhAqgbMICQA+NYg2PFbsYogD02ARWKu20CxW7MBWirMICkG/ySqI1WHK9C6W8GjiFEHkjYSGEcEXCQgjhioSFEMIVCQshhCsSFkIIVyQshBCuSFgIIVyRsBBCuFL8sDAUKhIsdilEgahYqNhFEHNU3LAwDMyGhAzhrgQKjPrqYpdCfAjFGxvi82IkYlj9SchNFq0YogBMA6O+Gjs5BhOyFMTpqihhoYI+jHgUq3eo7GsVGo0yTfB6nMlsK23ck9fErKvG6pelIE53RQqLANahwbKfzFdFgxiRkDMS1rYhFsbuHSp2sQpKhYLOl4LM8H7aK0pY2IMjhT2goQo+dF2jMaNhrO4BtNYoQFVHMRJV2APDBS1LMWmZX6RsFP9pSJ6pkB8VLvzTFuX1oictmAoKAHtoFOX3OnOFzidDoarC4Cu/6UlE6Sj7sCjWVPkq5D8y5duRnxnKWcB3vttpfF6MeLTs239EcZV/WBSJHklhBP0YwalFp5WzgLDOx9MABViWM5O4EHki9dZ80WD1DGE2VKOrws7PbBt7MA9rkNra+eOR7Bf5U35h8cH7dnP2Jf4Kwrad9T+VQlt2/iaWzeTQmWxRVi4vKq8J6ph31TSLV5YKUF5h4fc6jyqPbSnQYKeLuDSArQGd9xmodW6ystosTAMjFuHYa21oT+X1Yymg8gqLTA47UzmPJY+lxyqsVmHZMx5BK48fojLOKF9OPSyUQsXDKJ8P5TWdzlXS4ab47PzUKlQsjAr4UF4P9uAweqKEFnASBXXKLWIapwem3Z/ETqWdbsyibKlQADs5ijU0CvK0paKdevO5to+2vmdzKAmL8pabBBTk5FpXulMOC4Vybjs8Jjqbc3okirKlszmUz4POWRIWFW5OD+YPf4CwbDCMsm6A1lR2A7tzrb3O0xytK/q9qHRzC4tMDvw+tK2dcQllvDKtUmAc7lRViXKTR/qu6EmpXVSyuXX5m5xEeU2U1wSU684wgeZmmq+8kEBVYE6HPRnl8WAGA5gubo2Uabrb1jQxwgGUx4M62QAww8AM+DEDflx1rFAKwzP7e2cEwzRcfiHxhY0n3sUpnPPhMp70PA5v5zGn+oko8JjOlALHCQsjFKHxiouo6qifrZREly6hcfU5mD7pOHW6mtPXhLZs54Mej6JTE67mpai7Zj2r/uIOAhEf6f3v8fRt/4XUUAaUQbijjVBthJF3dpEZOdX+AorIkjPovOmjNK/5CJHWOqyxEfb//BG2fOeRDxRNEeroYOGt19J06QpiCxqw0ykOPPprtnzrZ1iTmlDnQto/vhqTLPv+5QlGDgwRbTmDc//yNoIRg50P/Yj3Ht8yrQS+RB1tn7iGBesvJn5GG4ayGNi8mZfu/yvGkxk81Qk6PrGOUHWAQ09vpPf1PfhbO1j5tS9Ss6iO7l89xta//jX21DB6X0Mrq77/AA3LmtG5NFvu/Tq7n9p+SuccWbKEBR+7GJUZY8/DT5DqHSVxxVpWfOUmfGaO7d/5AXs3bCPQ3MqC6y/DH1AceOxJhnb1Ell2Div/+A+I1gbZ8+N/5J0n3sCoiaG0QXxJKx47y9C2XVg553FtYMFCVn33furObMTOpHj5Sw+w7/ldTlENDwvv+APOvesGTBMGnv0Nz9z9/XKfyqQsqf959nrdYfvzeASTts/czPn33YLXP5VNWrPlrvvY++YQKx64iwXrzsXjNRjf8x4bP/91RnrczYEQWriYZXd9hgXrzsPj/0DuaYtNn7mD7rf6AAi0LmDZXZ+lff0FeIO+Gdu+dOe9pPyLWfXnXyA4VfNJ79nGxvt/wuqH/oRwtfMza7SfJ66/m9G+CcxYnEWfu4kzb72KYPXMW5Vdf/19dvxmH5d85z5qOmsBsCdG2PSFr7Pkj79Kw/ImZ0PbYvMd/5F9L+wlctZHWPWte6juSBzZT//jv+KZr/7Q3Tnf9kewcDUXfu338Yed80xtf5Xnv/E4lz10P4Go87PJgf288Kf/xMr/eheRWqfs2d59bPrK9zj/Lx+gqjnm7DI7zoZP30na38r5X/8j6pYvQClN31NPsvHe7xE66zxWf/seYs1VR4rR/bN/YtODP0UFwiy/726W3LIGw3CqWjqX5skrbyM5NP99c0yPn2C0dt73Kxx5vQH1VCU452t3s/Da8498WAC0nkTVtnDFP9xPTcfRixvqXMyiT1zCa//niRPu11tTyxlfvI0zb12H13+caq0y8FWF8MTiLPrDW1n6H9bjCx6vqm7QdP31NF5zJV7/0Sp6oH0Za3/wNbzRo7dNRjhKsK6G+NqLOPuumwjXRY/bZlO18nwu+9TniDVGjv7/QJRL/uYbeKJHZ7nWyiDc1kRr64Wcd99njvySHzaRTLo8Z5MFt99G88euxOM9eh6hpStZ+9AyvNGj+/UkWlnz3Xsxjhl85qtr47If/Nm0silvgPbbb6X5+msIHCmXonbdOs5/0EPT+stmvK8TySTBjkVc+M3/RP3ZbdPeH50bJZ2STnyno7zULIxgmJaPX8VZd95ErDk+43VtWeRSGXwzpoXX7Pgf3+LNH2+adb9mJMaCT32cZZ+/gXBtZNZtDrNTg7z9w9/QccvHiTZVnXBb59AaNy21OptmZP8gsYXNJ9/c5T4BxvYcINzROktTh2bgxS0EFi856Tmf6jHzQ9P/4mtEli8nEJ35ucrseYdnv/xthncfmvcjS80iv+Y/LDwBLv6bb9K2auEcPrOagWefYuM93yeXmf7tY1TVccWP/zu1i2c2oNm2hWG4azg7lW3d0toCzIL+jubjPArFzkzwxp9+k52PvTav+5WwyK95nwDBW99By5yCAkCRuPwqWi5omfFKfMV5JBZNDwo7Pc7en/2S3f++9aR7trMZDjzyK3Y+/OJcCjYrbVsMvvgir3/n4YL1PziVcy5Vhj9Iy3Wri10McYrmPSwmBw7Q924vWmu0thl6bStjg+Mu/7dG5yaY6E/NeGX0vXcZH0k7+53M0bvhOTZ89h5eevAnxFcsO/4etcXAi5vZ+Ll7eeGBHxFZduYcz2y61O73eOXeB3n6i/8Ns6EF40PWKrTWZAf76Xvz/dleBCtH77PuzrkwNFZygP7te2d5SaMns/T87pVZl4RxQvbN/BdRzKt5b+DUmTFe/ML9NF+xkol9e+jfuoeLfvRdIjVH2ycmDhygf9s+6i+9EH/I68xLiSa5ZSs7//5het4ZmLHfXNf7bPjsf6Zx1VJG3trGwNt7px6/Kca7BqCldfr2Q4N0Pf0CB594nu7n38K29NS2/bC8bnqZ0U43djfnZ1sc/Oef88q3f05u3FkHY/xg78ztnCF3ruexSL7xGpvv+99UXXkjted0onACxE6n2P+rp9j32AZ6X9+Fto9/zqdyHm5prRndtY/IonYM5fxbZ9P0bHiBHX/7M8KXXkdiWfuRo1qpEfb+8rfse3wDgwfSXPP4Q3jjhxtANcktr7Pj//6SgxslLE43+X90CkTPXslFf34HXpVm908fZdcjG7FyNrEVK1l042qyhw5y4N83Mby/f059q/2tHZz9pVuI1IUZffd9Dv3uFXpe3oGVmfm15q1t4ux7bifWFGNs1156nn+VtF3LFd/78vQnNrZF/6bNGI2dVC9qQGmb8X172f5Xf8/7T7w+rZzKF2LJXbfTsKKDiYNd9L/8Bt2vdXP1w98iEDzarqC1JrVzB8leTdPFSzBMRXagn/f/3y/Y9o9PQzyGHoeVD9xN08o2ep7eyPYfPMxY78yp+GY758lIJ5f/ry+gjrkH1JZFz9ObCCw5m1hrDdiTTHT14m9uxuNR08qWfHULWW/iyOPRdHcX7/7tT9j56Es0XXs1TRcsZPitbRx48iXSSae2aERruOCb91K3pJ5Dv93A9r97lPFjaoZN19/Aii/dSO7Qft754T9zcNO2vPWxkDaL/CpIWJQ808fy+7/CkpvXYCjN6Hu72PmjX7Dn315CGz6inc0oO8foni7sSffzRrTeeivn3fNpfBEf6YNd7P3lv/LOP/yGbNoivKAFb8Akta+L3PjUHBEeE7MujjU4Apk5rN7lCbDyG1+l82PnYWAxvG0H7/7dz9n35OsoX5BIRxPk0ozt62PRnZ9n+R9eg8drkNq7l90/+Rfe+8UGLDxEO5oxDM3YnoNY2dPnMaeERX5JWBymDPy1cQylyQyNYOfm55fEW12Fx+chNzLKpJuJY0wDs6HGmbtzLtPkGSaBRBywyQ4NnyDcFP5E3KndDI/MWgsrlKkO5R+ahEV+le6ooIAPoyoCk1ZhVvDSNpm+wXnfbW5omFOqI1g2k119c297sC3SfTPbfGbSZAZKYylF5TExaqtAa+ye0iiTmKl0547PTqL8XoxIgA/9qOE0M9+NlKVOT1oo08AI+CAgs3GVqtKtWdg21sE+px3Rzv/s2KJ4FDhrwioFdh6XTBAfSumGBUA+19oQpcXWKJlap6SV7m2IEKKkSFgIIVyRsPgADU6DqmmAz4MKuZz1qhC8ptMAWCrlERWltNssCkyFApjVUfSk5YzHMAxnnMN4HlY+P9WyhQOoaBiyOYhHsA/N/2NeIU5EahbH0ONp9EQGnc1i9zrP++3BkSKXyqGiIey+IazBYaez1nHm7hQiXyQsPsAaHEF5vRh1VZDLMeuwySLQmRwqGkL5fSift7IWQRYlYfawMIyK6wh1mALsviQYBnbS3VyghaCTzmAyIxrC6ku6miTZFTXVPiPESczaZmE21oDWWN1uug2XIa2xeoZKqx1Rg06OzXtPBCMRQwX9WAf65i+ARFmaNSzs5GhlL8NF5TxwsEfGUemsBIU4qVnDohRa/0WBZHPo7ByGw4uKIzerQghXJCyEEK5IWAghXJGwEEK4ImEhhHBFwkII4YqEhRDCldMsLBS+6tjxXzY9+KrCc9+9YRJbdgbxRU2ndHzD75923EBjE3UXLMU45t1Vpgd/oppwSwP++EnK6PHiiwXncALgiUYwvNMvq+HzEahPEG6pxxs+8UzuRjCEJ/DB7jcKX40zE7ioXOY19Yv+LK5Lb6S6Jxan+epLCEQUqUNJAGpWraLzoysYeHU7/uZWWq6+GMaTZIYnwPTS+nvrqVtczcD2/fjr62m49AJaLl3O0Fs7T9pBUXkDtN98LYll7VQ1xxjaPXDC42sN/oZGGi+7gAXXXU68LUz/G3uoufgi2tadS3z5GYxsfRMz0UjjFRfRtv4SYp3NhNuaabrsXJJb38bKaUIdnbSsu5DJoT6yY1nw+FnwyWuJN/kZ2tl9/AIbJomLz6dhZQcj7x1Aa/DVNXLm524gu/990iMZomcupnndJbSsPZ9IWwPRxZ00nttG75adgKLqI+fQvHo54/sOYOVszFg1i2+/ATMzyNihEZTXT/ycpbReexkt6y4ivedd0sOl22HPMDx4/aGTbyjmpPRSYkrzx64gGA9ipHrA9FB/+RpaVi9leMurVK+5jKYVLViGj7E3DYxAiLYbriGxpImux35L26dvIFbrZbQ3hc6ksCwIL1xE21UreP+nvyaTmtljsfGatVgHdpPxL8dMw9LP34CVmSQ12/FXr6b54jPJDScZ3LqDQy9lqao1aL7uamIJg/63D9JwdiNNn7yBQFDR/8pbvPPUc0xO5Ah2nknnVWdg1jTQcvlSEssasfAxtBnMcJQFn1xPdWcd+x95nfabf4/hzRtJ7pu5FELsIyuoXdqKL+SkYKhjIZ2fXIvHHsXyxjnrKzdiDfXS9+pb7Hv0AHbOombNGqprJoks6qTugrMJVvsxQ35A46trYOEtHyUYMziUtDnzi7fhD5uM7d5Lz4bNeK67HDPeTMvCRXQ981qljwaoSPNfswj4YPLDL9Az8u5ealYuZfCN92j66Fr8apSJMUWkvQUzl2TPE1upXlRLck+S9k9cSXr3TsxEHZG2JtK7drD70efwt7SjRwaJnrOC+uXNHPjXDUwcZ5Hm8T17GD44RGxxG9mBXrqfe53o4vbjHH+Evb9+lu5NW0l19VN36SqiLTWM79rF/idfxtfQhEGOwVffoOuZlxg90HdksZ+6NRcRa6sllIiS2ruXvjcPEmsMMtKbpePGKxh7azu+liYirY2k3tlG/7aDs5Y3c6gbo7qJyd6D+NsX03zRQvq37iLW2Ua4KU7Xvz3Fwee2MtE3jLY1KJPm9WsINSTwhz0k39rB2JCNN5fECtay4Orz6H/5bSKdbUQXNND/u80ceOIFBt9+HxWuoXnVWZimzcDrO8iMTDiF8HvBLp2h8lKzyK95X5HMbKnDOtj3ofdjhGMsu/Nm9OgQvb97hYFt+zAjUbwBg4n+YfwLFrHstrVMHOyme8NmRvYP4KutQeXSZIadQGi96Uaqm4P0v/wGva/swMq5/2Cf7PjHfrVGFraTOdR1ZKHkE+7X58PwKCanxt+Ely7njBtXMb5/P13PvMRYdxJ/XQKdHic7OnHCfbV86noS7VUk395B98at5LKaUH2cTP8Q1iwrqpnBANgW1tTSiLVXrqXl/HZGdu6i65lXyYxlCNYnyCWTTKaPnosZiRFOBBnZ1zPtvM3GBFbfUMnMrSErkuVXyYaFKH1GQw12f1LCokLM+9MQPY/VUq1wpo+r0Il4St48DmvX4Fxr05D2kBI17w2cVvfAvMwFocJBzKowOjeJ8njQmWzJzIcpHNbUPKUf+nr7vXhqq9C5STBMsG2nxmJLbJSSeQ+LeakDeD0YVWGs7n5nhijAqI6iqsLo4dR8HOH04vWUzFygx5qXa20ozNo41qGBI7czKhzASFRh9SUrZhKi00FJdsoyIkHsoaOzdSmcOSiN8Nw6Kp3W/F6MSPmetwr6sVMT09o9dCoNpomS28+SUpJhgVIz2j60rryZ/jRg1sTQ5TzlnVIzbjc0TLWHSFiUkpIMCzs1gRGPTPuZEQuj09kilag4jFgYDShVvr80eiLj1JyOqUWoqVXX5rOxXHx4pdmDM5NDZ3IYTQlIZ517dgV2b7LYJSsc03Bux4bHnHVCypVlYw+PYTYm0BMZ5/bDa0p7RQkqzbAA7OQYanQcfB5ITUC29Br48kUDZnXUWbeknG9BpuhUGmsiAz6vc74ZmUC4FJVsWChwGr0mKuvWA6aq4aaBPZ7GCM5fh7mSZmunFilKVsmGRUEZCm3rkqn2mjUxUApPUwIMw3k6IESRSVgAKhrG8Hux+4dLYmDUjJXgKuBWRJS+knwaUmh6eMxpZGuoRkWCxX9Eq/X0P0KUAAmLwzI5pxehx8RsqHHGKQghjpDbkGMdXnx4akDTfMzLIUS5OHnNwleBeTJpVebjO68pnSbFcR03LDSgYmHMhhpUTGYfKncq6MdsTGDUVBW7KKJEHTcszLo4yufFOtjvDOAK+ApZLlFARjyCqopgdfWDoVDR8h24JuZu1rBQVWFQYPUnwbaxepOYiSpp9CtHQT8qHMTucYaI2/3DGJGQfDmIGWYNCz2cQhkmKuT0HlSxEHrSKok+CGKeTWTQ6Swq5gzcU+GAMxLUksZdMd1xWy+t3iHMxhp0NAzZHFbPoLR9lSlrYBhPYwLt84BSTqcw6d8hPsBjodMoAjN6Itk2Vn8S5fOixyYkKMqYAqzeQVQ0jB4eK3ZxRIny7E4l/0SF4w+ahprZqmVlYAKQporKMJY+ra91xDRpL3Yhytj/B/IL7tRUCZUiAAAAAElFTkSuQmCC"}]}
