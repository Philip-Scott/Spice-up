{"current-slide":0, "aspect-ratio":-1, "slides": [{"background-color":"#ffffff", "background-pattern":"" , "items": [ {"x": -624,"y": 442,"w": 2791,"h": 472,"type":"text","text": "","text-data": "{title}","font": "raleway","color": "#000000","font-size": 42, "font-style":"regular", "justification": 1 }, {"x": -621,"y": 771,"w": 2768,"h": 315,"type":"text","text": "","text-data": "{subtitle}","font": "raleway","color": "#505050","font-size": 28, "font-style":"regular", "justification": 1 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAWwUlEQVR4nO3dd2AUdd7H8c9sSzabZBNCCr2DdEMnFAMJXUBEpEjzxK53iKLPqcehngUVO6iIcBKqSBM8CAcKCSEQRHqXQGgJIWWzKZtt83n+CIeGoj88CzzP9/UfZGfnNzO/fe9MNploEydO7BcXFzfLbrfXAKBBCCF+QKfTmZ2WljbBFBcX98nQoUNrGAyGP3pQQogbj0ayOslZBrvdXl1CIYS4Fk3TYLfbaxgglx5CiJ+nySmFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEELJTR8LknCVFqO03AP+YWPQ4XGXw+Vywef3X/eybnc5XK5y+Pz6bzTCSiuEz+uFy+WC2+MB+dvutf8cnzKF46P7/Sgvd8FVXg5d/+2PJkl4PW64XC54vT781K4gdTgL85CZeRIut+8nn9ftKkVxqesnt/dGmLfXy/RHD+CX+M8EP3V4JxYkzcOSZasR0f4urP3sdQQYtcseq8OvEyaj8Vddv9dVjPSUr7E5JRU7du1FTm4eXB4f7GGRGDz+L5j0p0EwadpVl/WUFSFt00ZsTk3Fzt37kZObh3KvjrAq0bhrwiT8eXRfGK6y7E/JO7Ebr3+4DJOmTkVM0A/bWrGvdJw4tAcbNm5E2tbtyMw6DYezFOZAGxq3isO0N/6BOhG2q45Vu8Y4SB+S3nsFlmb9MLxXe2iXLQcAJ/ZvR9K8eVi68l+oFT8Oa2ZNhfHi8/3nMY7cU/hmwwakbEnD/sPfI6/AAR1GRNesj6emvoY+7Rtd57iI3d8sw+q9JXj6sXEINFV+nO4rx3fpqfh60yZkfLsbZ87loMTlhi20Crr0uRsvP/8orD+eQyR0bylmT5+KV975FFm5Dtz5+OtY8u5Tlx1f4sLpo1g8fx7mL16G8vCW+Pe6JYgKNPzoqSq2OevgDiQlzcMXK7665ry9ISUnJ/NmoOs6dV3nhdPfc/5H05nQsSUNGmgwWWgygC0Sx9Hlq3gMdT+P7c3gtClPsnm9GFbrOJK+X2H9Pk8Z0zes5P2jBrNKcAAB0BwQzOat27JnQgITesYzJsxGS432PFfkrrSs113KlLVL+afht9NuNRMALdYQtri1HXsmJLBnj9sYGWJlQN3udJT7Ki1bmJ3Jd15+liNGjOL8tRnU9crjOrU/hW0bRhIwcOWewkv/fy5zP6e/MJmxTWoTAAEDq9dtxK7d45mYmMA2zRoSAF+an15pW/3ecqZ+tYgTxt3DR595hXklnkpf97lLOP3JEQTAbmP+Rv+PxpKTdZhzP3iN8e2aEgCNJguNBrDtoEfou3gMSx3n+fnc99n/tvY0GzUCYGiVaLbrGMeExETGd+tIC8DOI5+79Nz/ef7Mfen868SHeM+4+5lx9Pxlx8jPlOUzWcVmpK1uB55xeCrmjd/Lvds2cvIj41gr0k4ANJgC2LBpS8b36MmEhJ6sXz2CBlskNx92VFpfSd5JjkiMpcFoYefut9FmAtve/iDL/RXbUpyfzeVJH3FIrzhajBphNNNiAqMbdWW2S680bz+b+QZ7dmhO7eJ++fG8vdElJyfzpokFSY4bNoBVw4JpMJrZqEU7PvPS29zw1XxWMYHjpnxKZ0EOP/vgZfbp2oa2QAuNRhM1gB2HPckfH46yolwmzf6Yh04XKK97z6bljG/bjBaTgYEh4ewxYBhnfraUJ87ksMzlpl/XmZe5gw2rBrLtoEdY5q2YJAXnT3PhjGmMa92YZqOB1tAI9ho8ip8sWMGss+dZVu6mruvMPriZtcMC2GXEZHr8OnXdz7xzJ7ng41fZol4UjaaKbel615P0XtwYXde5P3UFW9QKr3jBNbiNTp/OglN7+djo21kl2ErNYGLD5u345JRpTN91kA5nCb0+P/0+N58b25MmWzV+fTCbJOlxFXNnylccP7QnLSYDjUYTYYli6uGcH/adI5t/vXcAjVpFfKYv3Ubd5+bqhe9x2IAerBJqo8FkYZNWHfn8q+9z3fLZtJs0PvL6YhblneWMF//CxjWjqAGsWr0eR93/F65ITmFufiHdHi91XeeWRdNogMZnPlxDnaTu9/LEkT187dkHGB1mpcloIgD+z/urL41L97m5/KMXGGGrCHGv8X+nV9d5OG05B8S3p9ViojnQxnZd+3DaB3N46PhplpS66PfrdBedZXzTaMY0T+D5sopQFxecZ/Ky2ezWuh4tQRF86cOFfHpML2rmEC7YuJubv1rIe0cNYY3IMBoMRtZq2JwPPzWVaVvXs67NyG73PMuyUgdXLpjJEYN7XZq3jVt24LMvv8v1q/5Zad6u+WIhz5yrHL8byU0XizoNbuHICRO5+ut0OsvcJHWueOcJAhrvHP0AW9avQYOmMbJWQ/752Vf5yZtP06SZ+eaSLSQrJt3e1NWMj21Eg8nC1xekKK/7o+fGs2pMXT44+SXuOnySPn/ldwPd7+aU8b0ImPnhl+ncuHoJHxx9J2vHRBAAw6Pq8PFnX+Peo6fo1y9b1ufipGFdaDAFc+66DCavWMD7RgxizaiKCETXbs3Jj4+lAQa++M+vqZP0e91cO/8txoRaaTKZCGh8+NX5zNq/hYlt61IzWhjX6w4uXZtCR0n5ZVuj80jKIgabwG53P8F9uzP45gtPs0OrJhWRMNs48sGn2bZOCOu2H8y8Ml/Fu2PWft4VH0uj0UiDBobV78zj53I4c+pDtJpBe1RNjnloMtduzmCxy0NSZ9I/7ieMFg4fez9vqR1NTdNYq0lrvvHRfJ4+X8DLdgXL8k+wS6OqDK3Vhtv3HeD8We9wYGIXhgUHEpqBt3YZzLGDulKzRvGbwxUvLk9ZEac/cy+DzCaajAZCC+Ci1GPc8uWnrB9joyUwhMMnTOLmHftZ7q18jqnrfia98hANmpGT3lrIjJR1fOrhcWxcpzoNGhhoq845a7Zx/9dJDLUYaI+pz3atGtNi1Gix2dlr6HguWfM184pKSercteoDGjQw4Y4x7BrbhEYNDKlajSMmTORXm7ZfmrdLXn/0h3nboAaNRhM3p6Qqz8ff200Xi8JiV6V/675S3tO9ycVTbLBFXB9+PH85cxxl1HWdrz0ygIHhdbnvfDlLC85wymOjGBpgYkhUfc5YlEy3z3+NNV3JU17KgqLia3695PReNqpiJjQLw0KCCIBhMXU56r4/c9GyL5mZfe2zmKLj6awZaqRmCKA92EoAjKjRgGMfnMQlK1Yz88wZju7RjLZabZld5meZI5vPPzSMgUaNTTr15wPDEqlZgjjmTxMYbbfSGlaT7y5YT+/lr8RL/HxxfA8CYEiInUYN1MxWxiUO4psz5jA1Yw8zVr1HA8C/z91IXfdx67+S2LRGFVpsEXzyb88z0gK27DaAfeNaUIOBPe9+jJnZRZcdn2IOblPr0vGJvW0gP138JXOdrmuMi9y59A1qAAOswQy0mAjNwPotOvDJv73GNeu/4enM3WxSNZBxd09iuU9n9rGdvKtHLAEDB45/nPEtajMgugnvv2cgg0wG1mjahf/ecazi8vQqfOVFTGxgJWCkPTSEAGi1R3LwiPv46YKl3Hv0FEny37Oeu3QpF9u1D6e9P5vfHsisvL26j1PGJVza3pq3tOX0j+fx+3OVj73uK+GwTvUrzdu5y5JZWu695n75o910sbicz5nFzk1jeEv7npy/JoVur+/S5YbuLWTPhhGsHzeEn814lY2qh9NotrLfqEd59FzhNSfPLx5LWQH/9tho9u4/mM+99AY3pn3H0nKP0nq8Jbmc/MBw9r19CKe8PJ2btu9lmfuHZU9++yXDAwwcOWkav5j7Lm+tH0OjOYjDH53KvFIP33lqGAFQM1rYtf8Ibj146mfWq3PLqllMTEjgnx5+gp8tXsUzFxz0+f3UdVL3lvLB/rG0VW/FtRuS+eg9/Rlg1Fi7eWf+a9th5mWmMdpacSkQVfsWvvDBQrq8V4bXW3iUrepWZasufbl43VZ6fH7+3N64kLmDwwb25pARY/nWjDncczSLXq/v0hnIl+8/RcDIN5P+xXdfeILV7EG02qP5wodf0FWWzyGdGxEAA0MiOPLhZ3kqr/gn16n7PfzopceZ2Kc/J/7PVK5at5lFpeVXnP25Swu58vNF/PbgCfp8/ivOiEhS95RyZM9GrN20Pd/9bCWdLs9V1+0tymTbRlFXnbc3qps+FtR1Flw4T2fZ5afZpPv8TsbYLRWnzEYzW8X15ufrt11xGnoz2LrsdRoABtlsNBhNbNq+BxddfPGRpMuZz/QtKdx3+DjLPf/99vmKz/G25hE0mi20BpgYElGNE55+lecKSipi4vfx+MFd3JK+g7kFzqu+cEiSus683ByWuNzXeMD10jntz/0JaAwODqI50MYed4xl+oGTF7+xrTM/+yQ3b05h5pmcKy4Vf3O6TmfBBRY6y669Ty4+Lj8356rz9kaVnJxMLTk5mb179/5dPnn5PdFXhtnvvImj+T50S+iDhG4dYQu4KT8phsuRjVkzP8TpIh1xPXohsXtnhAZZfrP1kX5sS/4Cn69LR81GrdC/fz/cUrcarvPT3N9E9rGdmDl7IWiLQu9+A9Apthksppv+x4VueOvXr8f/2VgIIX4969evv/l/glMI8fuQWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSixsM6UdhoQP+67y7tdfjvrQMqcPpKITHV/lu4brfB0dhARxFxdB/47t6V0LC43YhPz8fpS73L3oKv9cD72XbQ92P4iIHCn5if/14v4j/zs35O9u/M93vReaRQ/AEVEHTBjWhAcg7dRBzFq3FfROfQLjRj5yzWdi5ez/ax/dHjN0CkigrLsShfbvgNEajR6cW+Onf8CZKC7Ixb86n2HkwEyMnvohOdaw4dCQTDVvcirAgC6h78c3KJOTYmmFUn07wecpx+uQxpKVsxrZvD2LU48+ibV0bli2Yi80Z+9F12MO4u3tTHD2wG1vTt+PEmVxAA0qdTnQd8iCG97oV1H04dfwoivxBaHlLXWgAHDnH8cknCzH6qedQzXrt9xN3aREOHTqKag2bITrMBtKPnRtXYntuAB4dOQCOvGzszNiGb3ftRYHTBWg6nGUanp7yAupFWuEpc+LQ4SOIrHMLqkeEgNRxIH0dNhwpx8R774Tu8yLnbBa2b01FaloGOg6cgKE9muPk94ewJXULjp44Cx2Au6wYddoNxF/G9IWmAX6vG6dPHsPW1BSk79iHYQ/9Fd1b1/5V58T/RxKLn0HqWL90NlZs3IGQht3w+tPjcepQBt5+ewZYowOKju3A9Lmfw6MBeYVuxPa8He4yB5bPmYuMzDPwlOSjZZ/70EP348TBb5F+vAgjBvW64lb/Lkc23pr2Nuq0ag3L9xdQeGwb/v7JJuQWFmDC8+8hrl4Q1iycjYVrUnHv5M5Y9c+Z2LL/OALt0ejSORa2vYdRcuEUXpu3GNFN2iM4IBCGkjOY8kwSgms2RHx8AoaOro+wIOCtl15AcJABO7ZswIaN3+D02fPQo1tj5ouPIfv4Hrz79vvItdSHL/sglh/Kx+D+t+HyO9XT68Rbr7yEo6ezMfDBKbijUz18vSIJcz9fh15jJyL5i7lYk7ofLdt3wsDh41CnZnUUn9mD1z5eA19JDr5K2YqNmzPgKMpH4tjJGBHfDFvXLcWspJXoMuxhbF2zGF9u/hYICEGHzl0QFbITfm8Rpk+dAocpDD0SE9D3zkaICLNhycyX4Q614cB3W7F5UwpOZl9AQGgkunRui+A9+1FWdA6r1h5F394JN8ct929QxjFjxkxt0KDBHz2OG5YGICyqJgoy96F1977I3rMBc1ekINIeiDJXGTK+O4IhYx5AYptq+N4RgGbhbrz37gyYa7XEAxPGImtPBjok9Ebal/OwYtMBJPTug2oRoVf9uxe1m8YipDwTKbuOw2aPRM+urXDiPNGvc33888P3kGsIQ8G5PBTlHEGZrQ7GjR+PIbf3RhgcWLZyHbKLXEi8cyTa1CDWfPMdzIHB6D9kFEYO7Y+6NWMQZA1AQdYBLFixHudzzqKcVrTr1A0293k07tATzu/TMWvxOlQND4HLXY5t23ehY49eqB0dfsVZkWYwoXaNqth/OBv9Etpjxdz3ccBhhKegAK6iszjnCsbEJychvtOtiIwIh8VsQtpXn2P7wRPIyjqN8Or10L1zW5zKyka/Pt2wOmkGdpx2A6VOuJw5OFZgxOixYzF86CA0qWXDwnmLceqCA5163Y4J996DJvVqIthmha/0AubMno8LhXkoKPGhZWw7JPYdiDsH9kGEuQRfLF+L7IIStGrbAfVqRF7332MRFY4fPy43v1FBbyEmPTwJfls4GrbsgNEjhsCdexyHzzrRpm0s7EEWbF81BzNWbEPdxs0wfORINK0bDV/pBUx+bCIQUROd4vthUO9uP3u3Lt3vg9evw2I2Y/eGz/H2oo2Iia6GvkOGo3ubhtixJQUhNRqjaYNaMBoqJn5pYTaOnClGy2YNYTYaQN0Pj9cPs8V8xYuDug6PxwODyVzxh5f0Erz41GTk+gNRv2ksRo+6CwbnWez9Pgex7dsj3BZwzT/ok7VnE/7+dhKqRkajW78hGHDbrdiXkQ6/LQa3Nm8Ik7HyJYzf54XXr8NsNsNoMODc4XQ89+onqBIZhS597sCA+LY4tnsHSk3haNOqCcwXl9c9xdix5zhatW6BQLOp0h27SMLjccNgMMFkMlYaq6voPA6eLESrFo1hMhhuiDt93azkTlmqSDgK8uA3BiDcHnLVdyePqwSOEjfCq4RfmuTU/SjIz4clKBTBQYHXPVl9HhfyC50IDasCa4D519iSK5FwOgrgoRFVwu3X9c6r+zzIyy9EUGgYgq0B171q3edFfkEBAoPtCAkKvO7lxe9n/fr18j0LJZqGsIjIn3yIxRqMKGtw5cUMRkRERv3i1ZosVkRHW3/x8ko0DaHhEb9oUYPJgqjo6F+8aoPJjMioX768+H3JR6dCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUSCyGEEomFEEKJxEIIoURiIYRQIrEQQiiRWAghlEgshBBKJBZCCCUGAPyjByGEuOHR4HQ6c0jphRDi6kjC6XRmm9LS0u4jOctut9cAoP3RAxNC3FDodDqz09LSJvwvh2e7syBupfQAAAAASUVORK5CYII="}]}
