{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(to bottom, #164f86 0%, #5e337b 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/black-linen.png" , "items": [ {"x": 408,"y": 723,"w": 715,"h": 297,"type":"text","text": "Subtitle","font": "open sans","color": "#51a7fe","font-size": 21, "font-style":"light italic", "justification": 1 }, {"x": 49,"y": 514,"w": 1425,"h": 377,"type":"text","text": "Amazing Hipster","font": "raleway","color": "#ffffff","font-size": 28, "font-style":"regular", "justification": 1 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nHS9e7yuV1Ue+oz5fmvtnYTciCAIaqhgEBFBDQJyKQUNCEQFBY8FRQUqyNGqlWptT0u1p/rr8fysVvBXRKEqxSoGbEVABAEREEEEREHlIiE2QriEJHvvtb53jvPHGM8zxru2Z2nYa33fe5lzzHF5xmWOaZ9zr4c8d5y67NkY4xBwwAH4BMYCAA6fBhvwdQ+zAYfDbLj7ambD8zuz5cDjvuGY0wAHbIn7AbjPuB4OwBD/In8HHCsMS15nDhhgMPfpBrN8VtxsBrij/RvjgQEwhxnc92YY8LkCY8BggI2432e81wz83TFhtjjc6/k52Bhbzj3Hm/c7fJo+t8H78sdhY+dzHplhiXdovjOfwucOd6xmGPmcGeTPa2pMfv573JPeQTf31ZJ+bm7x3ViSViPG7BNmxr8B2Pl0bfOI64I2PvdaNzMrmsGc66hnjAHM9QTt+0+sg/sqGrrvY85Jgfqd9DNgDPg8htkO4tsgOOCr9TUK3iA1k57BJwY4ghY7wGe+Y3DpySOW14vPfE7YWMTHNhb3uVryEdwdpnW0Wjeg5goL/pprPqO9V/8iaR9r6pgYdgD3ueHfxh+WY/MQ32k2Yu3c3M2HYeS4jNesZlayE+uZ9PMJGI7mbTf/vN3xfo/9xNHBZVdgLPA580uDjZgwfAVsAdbjWt9lFwwwllAg+6P4jAQC4HMPW3bwdS2GCQUU98w13xXX6/u5j89sbAkWVA6iFAPrMz8+B1t2EjSfa8xh3accWMzDDFj3Gi98TR5eYbvD/CwENcYzY2FCMGo8Y8TwUhlpHl3QfAJjF3PignJOJ4TGlgP4eixBMBvxN58bTAP4DKZKGhosxkfamFE4tZbx3QJgpsI/QU/Oeexq7BzrXGFjl5fPej7vl8BQoa25NEuMbzlI5XLyJ54ffDaBOfPvXcx7jO24UiHEc/fx3nXf3i/BAtYj0REw+HqstdNajqbQ2jx8f5xCy/UK5RiKIX/P59iyKx4eKSPuwO4QmLFO3nmBPDj3erboKFngWqVhAGCj0TCEXHPw9TjGkWPT+oxdrgUNxRQQsOUwFO1Y4g2bNT/BF/meU8ef+tQOhkN3h80VBk9Nng/lovqEmwWjeWj3E2Jc1+ZLQmlYEzDTs8LSJ0NzgMtBWphgfBsWDKjFoHDupXRyZqEMdofxrBGKLJTDrpSEz3gHyBxkwBznWOJ7KQvENXZc86Rlh+W1s5hazNcUoFswP5Eav3Ok5ekWIa6tazwZerT3NmU5Z0MzOd8co3fm5II3y2a8bq7JaMmWvoYIe1PoKdTuXvchv8cs2rRf3IrJAPLCBgmdGBsFM64j88McvnqN3ZCGbFeKjTzE3+HAcohCx41bbQSPkz/HSCWFWsdd8kJMoJTzWFJZJb+kkaGi2AieDWDk+ywtvydPULl5vhMeBgkWxnXu4x1cc9LI8l2TY6VyFUqIcfvM2XoalD3MY84dnZL3LJ9P4xrILhV+yjviVYc7TIeNmQsVTBgLMLcPWdcwHgCw7mMw0wHsSzu754M9oFYKBgypZJayxoJnA8CMz1JY4z4rBqQFBVKgnO5QLNAkUQ0mRe7Aki+ftIhpWW3APBYI9Dbc614u0FwTXW1RjN7jon3CyuYemNW9eb1PDyZyh/kEbFfMOtek276g9lwBWyGrHRMrq+QTMAfWhM9kXEdDQ2nd6AFS6SQzxJqtpZxoJHwkvQyYFuONAcTzsU8UP9PK5u/kFyAs2wYqjy3RKFwN0ZblpaIhXVHXY8b6WbqXDjmIzuc19pFHlZqQSi/WO0ykzWYoZ4xXenrOdBdR68UfK16AW9LPpNx89UQYidgn+W6mELexzBn/ro1u7rnGIX8MBxAllFFYta7YHwNLjo1j9uT9GbzgOSc+w2qywGwuFA0iDDsbS9PSBlvS+pAhzWCW/i61oo1QGE2rW8JcEH5iCQFPJjerv80sCCbYlcqJC8lrqL1Hvmeusnqx0HmPWXOxqUWTSwiB3BNZz9S+S4QcgIS2SMbXDXxcE8yyhuV3NqbHLJdgEF2sOabZBIWci7L2qdED8tMNbIoh14RRjKDRLhg80YEl44dFK8Esy0h6lKU3W+DLkIWh+wBAFj7oazXORKExzuQFpDXV+w0OjsOSjKmciVITAbpQBUnTlUpDXz7TrYGUjDMe5WnwNvQtS1prWXwSyzZ1eTpGzQjti1chtVIPorIEYN55gYYwURmVsZUbVDyx5QPKmzuRd657IlcbS8rIKF7QuqWS3B2m4ofoHuMz2EhFoPd1ZBbyPXYHhXwbfQLXMNgFL212MsAli+PBWNaII//KxFzgtclgvM5spGKx/J3BxyXlYoFpcTojBPxUgJHXNvgakJGfmYTZYDLMEpJ0aywRR/+82MPb5zWusK6NCfXofBevdcDGgUaCpIUgIFB0z9+NAihamf4DZ2WNLrlW9XxNdOvmzHXzzD43PYeMzfE2xKix+gTQrKuYic8shar32Ij7kwE1RoPiXqJxU56aP8dD9wyBgmKtiq5UQiZLi1LaEZaUVabl1GcaUPJRdydPGIRNvCNV9EYp9edoHgh+pfvLOTaXWusKF+/3daXiLXeyDHGMb21jKWhV93HJ1npm8mk8L/VArnnEMF3X7DAdsBWeboegNv38dR9azWcG3JIB5x6eGsoV/EzblpoUS8Y4VgfWY7jHAvs64/6WEZCvPtewNJYCTLeI7g4cwBLMMCyFgApvB98fg26NB/aHDy5qMhADdGYRgKXCkHHLCHmH0wlT47r8nPBZSAYbKxi3HoFxnoDpnAeaq7amjM3GqBFxh5iZqMIz6DgyjhAIzNeZvvNQQNWbINuICLp7BlFznX09QsWihu4p3p/AOMjP8nmkGRA84F48kAFqb8rbGSR11xyFVNd90mTCJWxBcw/ORvpVcQ1jFysyiH64DegSHZ4MxM4VAY5yoRhKmKH8AsmtcZ0yR3TD6BbErb7uQSUoi8wg7QYtlCEI2B/rYhkvim/okgNwBilDCTrjC6kA3PO9K8hsQScmdkivuS8kx/eIFhO228HnVPCf8wv0WMF8F80n4NN2GJZZhLIIcTWDbAFhg7GXZuWXIJLFtaExTwgYEvrDgFEWMx5fEX0MpFvhpQAtiSeak6DNHaD1kBA3wdf1KyAitChziyqXcFNQmt+5HuWAimExPYOleU8LHCVHxtzp2qUilGtgmX1pCCLmne5UMpkNi+cRKXFhGWSztBrT4QNxvZloGz40USCRxq7WWAyf/utYQkdTIGfSiPeTPcZSynGkEOV1zoCgGTAOgnSjr23Mpaw2U7g9q5E8Il6M/2lTqXVUliAVBtdW9xKBbR6G0hZU2LPePLNMgBZaCmAFA56RxU+j6Chl1fmLQT5HjoFrmXyxcWu98UJ8bnmdkFpmFbcxEK75UkptUtZyXHKJJxyj3s2gO4P1XPcNMszrffgO0w3rHpUeW8W8yPsigFNSXMEPj4eNXcoTJ5kcQviT1wnypD8VtMiUFOH7mpp6ZmDFMs/Od45dWQFaZSA+J6HN8m+DMwrNcYtBl2QAWoEFzOcbNVaOzwUnUyg5LxDyJhN2P5DBIktNaIGG3HOe1q+DnmFjVwJKzU8FSOUsIcgx8t4MBDqtF8eVf1PpgP6yN/lyj+DbDEsuYfFItdFiM3OhILBqEpDpQsLsmpuukUA1eJ9z8vW4GRri4lTybulD5xqRdpiwwQwXlTb9/FE0yncotkVjwOzTFvBrHQfpNXZJvyVo4xnHM6DqQBhnOhETQPC7xk1eowKzUvyhEIkSPDN2jU9k4NI1syURHACv4H7o5ZC74AWIFwzIvzOoaiPQNQ27k/7MTM50/4GdhQkTM+hnJRyiZkUQzBHQJjMLymRIOy8NPiFhHpEAmWoNCClrkszESDMXfs6MDTT/ca7xZFpijncTVDIRnMwdvFfpSwrDRoGotiSi8RFYGi14ZVoEBeZUoGRaDM7ffcKcQrOWImUGgSiku2BIjT4Zj6DQ5DqoHoXCMbWooJLTd1REnmlCr3nQdZprWROLd1U8JMe17pN+NQ7NMyE1DYwzg9LjGmj1FCfjYQ0eI1ENlbNiScaVpmAAWDJewbqcXBunkHimhceArUWPsM5IAQY2NQsce4uheCJJW5hO7QqtODBqHqY+lwsmt4vrE2urORJ1AAByTJIDuss1d2fsEBZuhKf7Cdd6bGVtD9iu3kED0GivezNASl4oek74nDbCJaIAmR4mAafWZhxCEJGM2JkC6AzKwitLra5nS0gJO0MRGX3FbinSigQfjxonmdBaQNG6hWhjEZHImLkGVKVtzMFA6YeL6Jnt2SyEF+xLOhgVRLJRBRM7qqHiataCykZ0QqM/TvzdPp+znqhgJjQnKiaQEXgdHI7ZaF2RbyOU5ni1vrw2FH1lRDovoM0HNV54+OJN+PVsQfdGG/7vifiPPmtzjqBg5SvED2nolPLtwtLpoh8vy0/+5FpSKbcU5HnPmDOR1VKfixcg3hSfCuVxNjLr6NkqofNZ69CD4pqT1g3n/6RLE1815ZXyJSW+kQW0Zw4YzZ7cChYzIa15J5zpCY3I9W9fZv5IA1JxUDkYB2L6U1C7308tLwhWTCilID4r5CGBFtFp6f/hFGaPSHdBk4KbjZg5pn8orRnDqLiI7reeMiMpJyee/58Ii+9OmlQKdJ7HWkWAphjQ0VJ+32/saOP/V3CCjlE8bltBs4TgevVWmVj+btbWli/fGAwG0jjnrYKxvkaks21MAYK3msVmXQdamrIZuFIG8bk3oRaZMubjG+XS1lg8xCG0OEkWSCkL1dwt0mMj5P2nK8SmUEXPjAMZKvC4WeduSChfkt0yrp12vE/xwm4IaQjodcwVOy3W2NHdS55ogTCldOIlcY1XECUHueHJmgUY1KJNiwIXSxQ9W0Vmt5Qjo84Qs3gvOXfPmo59jLWVXcf4MrDp4gIwVqGoeypIZk16EDVGXbX/GyipObFasgT9PMjYrcTch499QmCtpX71rhOMvQ3skZ4uCgsdkKZECoqjZExjUPhnWTjbyZWgqIICQ8RHpWEjou+su+CIcp6+Uei1/kWLbZaGP1VD0n98cz/mjDJ9ojoWgDF46BFvwZyq55EAia5pGK3z41aJOYPWynKswDhV99H1q9k3Y+cRYASgAKhFQLvQRSAtxls0a7n7EI2i9iZdpMEYBV0Y1m/k+jZUoNjSzNBArlaX4zEW+DS4RQxHoIADGlkLM3awZcEushETPo/J40mw/Jnpnyr9tQK7BslBgc+/12ZRQWXa4BWjuRmNLkjXoK+Yv7kqZuXjd3u1EQYyIAXFNoyMTYwETcAYaa84hgQFBqV4W7CTFkWBw6YUQiFlhsEMNmNuroAV58J354I4i6oocFRaJvps6js6wutojcJDa6HHNXRGuk6HZ0rZJ1OH9KXjuuBbKjbuEyq6bdwPunuDAlK1EjXm5tYhDdV6LLqqDgCAsnIGrZs21rWALXTt3PINDEwDVr0Bg9sDhk6Tul5/M8vQ56egZLPsGQAHvMrIhYhQLvYm6Gpaunh1liEwWM/rOSYaFyvFrTUGco4AkaylAfMeQpArPTH35IHZjENNiUjf12NgzkAWZrkhjNYGO6VbHPsgqy1Ru0443OIEwxrhTliLTB+AWo2wZhjrCHhdMJKldY6cv2uRCKe0RwHIgKCHMIZWgCk4lM+T6zSzwhCwVpTCzXJRbtvKysGMwtwEA0P5TRkTQcLRhTBLeUH7n+OYTt4Bo9gxr0ULfl7BVactmZd0pqAaWhCOzMn0HjexLWKkoJ1lgmuIVjDLIimir+aCWqI4FKMzQO3MdEmJZuyAe3GQz89rpDgUZyGTUinIasVlYySvz4rTeAYm3WUBk0KoNGTc45N8wAuyhJ5rSUNB3ugFe45cRTQDmdBd+0OC78QL5KFZ9To0tirDT153CTF12JJzmKVgOIfcL1Wl2cE7tsS2gSrCS8SVSot7jrQxlPygjXCtYhNhVGJbhIGK3dywU8BwjAhh0OJzQbkDT5ty8kUq7bW28Qfl/68Fv+TjdrVlW21ZsJAC4PV8Ck9PlfJHlnOCm2x6MRORUjEsX0+rZPV9zrkWMT7jRjsoBqFB5iWj3V6oqvxHz81V9cx+u6wF2vMz5VoWqc0XVAZJdh+B7Mi4eU+sfTKN0pccc/mz5p2+VIS7CuA2puF8qgpzlICjrT8qhany+1lr59g+hz65MiugIm7/IZ9HxZB8ov0S2Aalld3Q3E7wTOM9KjgpcW3mIo+2kXc3qvGUfmxI6WxiPnApAo2V/GBdQZI32/MGeYJz2cdt06HCRTLEGDL2ljuYJ+t6DOBmSypvKZfN74wbZSxmHmCnDybaxB3O3LJ8plYlN/cthZeR8cW2AUpfgwnp4wE1QKAtoNfASkUVI7HegiTkVuENoxngCwR5R9uKrOAsQrPPFWB9PJBwON0P7dozDAaG0kIWDXJsmRbjeAtQxT3hrlB/tABqWnj6yiYNifqFY+fa0K2QssrKU59NeLzm7dvn+NrqH5oVRVeAfD9/n1WVi02KN9dI/JD3UVjXY7BAT+5ZWwvGHiTE3t9PPUwEZhpTubaZAYsFLeuZippogO6cwaodARdqOZBy7nteYMhiO2xdjKW2EMBG7k+hsHVFH2MyIGImYowYu/7OYsPBdUjUGSRMxaW1B1I4Y70dVYjGdYdLgSqWQ9Q3Z3gHPsPlTPQcKH5NsgQa2RrVoXFF7GWPnU83t1m+DstN5z6G4ROYfNjQgoVSb0zZFrx8n4RQ3f/yiSrY6RCV7NrcjAwk2bTwgc97D0qbMjgl9JGMyp2j/T3umqdKXZmtaTQI4lYfAVqqbTmx5aIUb3V/0pWqghCKNtP1DFH3FzscHKZ3lGVsz+/rQcWTQu0Sfmtp3irIcsyKk/R1TNenmrKwchcAGwp57jRFzqtDJY0PZekp7NqHk9e2YOymhsEWRHkzpJzkclrjhTUVotBnUz4zAq5Ct4ascch+DzRGJ9aUm/Gk+PfHUZHE77JEXUpXCmFWbGTO2JWeSnVjbHPebsk/zq0EVZGs9gFymYJm2r0td4kIalRMiuT1iLfJFfakbbrXaLEo1JtTORcq506QnQ1gLIsEx1KzCpplxeH0iTFyv302tWGhCnc+0jqbW2wfthHMPpawo31RELES79bNLKoFQWi1wHYZG+mEoWsE+oS7hh4WYNLntjBwSy9TZ4Q3EYoswZLXQcrNhsHtICzXcpCLm6nNsavr0tcvik8poBhbMrqzkjAW1g5ik5ki5bonKwF3h7JGzD5VMZzDfWSwOFEX58fAmQK60DO7OxdeaO0yLUHN4C13q8LAfgw2BgJ7LUIOpqBvKp4x2rsNlUJk9iXTcZ6/C/JmMDldXO6mjXGZ5gf3yoTRKABQ9y/9np+zwM6zVJvxjrFoT1S1PqgAp+5fwgWL3blBP/XqyCn2IK3ZSNkYgOUeJt8FOdizAgeSGXD9FHsx2O4g+CTRMpG0j4wVsbEPTHxL1DdRsabhC2A7GZ0Y264MuhCen+c2GXlhDODYsYNbQA36RLIOXKUKREZRCjJw5vlv/m1r3lMWg01QkJDZlc0IpnTrNRE5yOnbWnZ20kOzJp4ZBMLgmfc1ft/EIdTfwOJ5+QxpVVk9WiTCMSIgRERYig5FYKbpSCul1GYy39qqFPNZxnk01KVxIBRxWiNZLrkegVYoNPpsrtX0pfvRUlzbuAznzzXd+vUuIe4ggDxgCfM7YwXSLCQYijUFzqnUGU8qH56GoSx0rkOPTxm3sw/4mnAcJl7xWS5frG+iF/GRy+qqPNryfiEKL34QnQr9Uvk4MwcqTycvMfjqAF1ySwu+JjK37AvD8YCoNf7HvcWnfOYSZf+LNCROI0YBVdXvAlU3zzUUZPLjEAIlLWgcWlwGUAC+DFIhXjNDOLIMcnYBIiGmy7pwx2jfFm5jSVnMgJwxtwsJoXaablJaPWbRov3WmDoViDZc0UfUYjIQ652ft5DY8hP32MwGpJUCqvsTyiduAULkGwIVp+UQE2WqTFmQrTXSohfkKctnLR0LcjmVomuDTxX3WHuW53xH0cqtbQbE5r3BSIZOj7BYgGIecL3HEYV5QoGai2mt3Ca0OZxjFKrsa88VYaGZCY3IfdTcmpBK8mtVmUnosYRCAO06zuXEu6XkLbtHMR5FPu78oPETtZaRqO30zBZCaKLaRkYspOjO+RKG8N1cXw62rwPn1WInlgmINE5mA9MZ+yqEBVswmL63IdmMn22wWzuNrd6hYKqvibTCcIwqeU4L4emXiSGT4GJEapumaTcLVsTQ7/qZZbGsaVHFMsj8LQBgKGtNglgjshcsj3u32RLBvM6QXEMxULKyMbVL65WvZSHTZi5JM1/bO3uWQOKhv7krVIqISnozrn/gXUIzDqAgvz4zzrOskujJPoyykhUrcTbrQeylQGvoQ9+1rBDH0+ZIOsym+FvMQ9faQKHWLhxoCrHNtUFkT9pK0eZ2fmE5a3URG7q5nkMrXP54G3vS3DXWUmbM7LiKn4rvSrXV+9wnVNNQC48K9tb9vVaH9FAQWiw02pxSIVMxORJtleIqS5Hrx98ZvPQpepK/XXxCRJprfjIZAWDH6VTulkxOYQw9l2ym6ZNcpdHqu83CJ7zbMAUtFRclrVVY37Usu2ICoxGMkDM1+8i3UvMzp4yY7GDxy2zVm3137Ea4kWMNVbmp86dgW3U6j+dioxxFt7QC1gWFNE4LLLTjWfNA6N3HJGtBGsfzrNMRA8B64t1IARglXKlIZGNUGESklP0XG34q5mwwtrlMopkYnmOr+AGVLt9/slu5NbrEDZ6KItEK/fasGQgeYRYkLOMYS7m5jo1FZJu8yHDRv28I0GdzWVAW3YNnDKPo0Cw7dxITrUV2g9WVsxSJUWFQqGn1DUDsZFU3ra4UYOni5mooJZ6xkI46ktLkUWWbtK4c9xB/x08z9kL6LTaUsmvuvuNktvXuqcl7ARCbv6CYRpqIEVpGWT0amVhqsmqqQgaxYvS5wgctYdNsyXCKIqtfIODefGufrex7ga9HekZFq9Pn9doFOJbDzZxba/zMoEzMuUfPu7N+I8YfQiWL1Ldhg6RZw93I7fRqhEolpHet1MvJZNnBWtAfmVrbgRkSb9Y/bmQ2oaxxY6EadzJ6pNSydoJMM1pPUO9rzSg7FU6rh5CA5rVzboNybY/RxnrxuY5QDqqSFAuKJzzXOvz/GMvcHxV/ABH7OZEKrpha7UyFRbWysf9G7oeSlXXHpJsCwMGNc3sJnQoY/RhUdj5XMFA9Z8S3XAglgpriYYuMm0uoT6AA8qSA9oms2QqoBaPcueSlkbzcninZYtUwOjtE2QARRmRy2r3VEMl28fLcLm6thwELNzKIF5mSCvBo4LBMZ82We3ctdgwvhXWh5kp2cAoZNXlTIrQ07BTdeyDIovX7EnVk1H+Mg2YlU9vCEl10FABZSX4/cw+JaGAZ/Yfr+fxu455xrs1Ni2yDp+DULlRPxMb5nLTe6ZWCZ1oICgMSCvYjiD4ZDnCPS7oFzK64uWiQUpH/5NpSMeyPSzGw50jnLO63YSUrKkbFbtayqCuvAaq+ZREi2qZa0awueQNV3p/8UoqN8+4C0fgh3auKkSy6zvIa/kvAZRs/PpGA3PDMftgA2FqBwiZUa8lG6b63s2ao0NUUaNLiswI2f+Y8nxckZ2QNqzEzUDoainVknDGVyGQ2Jk2br4Avdb8UCyp24R61HGnw2Ptltyw77G3XtFQGcKwEO+iV9epjp5ulMc0yEDQyvZraceRmsDEwkGcbaE9ICgOKKFFBl9rPCMeWWuTWKr/6AYSCYAN0RXGBvLcIqb0fgpotvWeccz2jp+UsGZT5erMBSPklbGZaN3Wn3AhbspGK17g1zbEZo7oz5XtH0rWsAAusEEIRE4V1AViK2TSXvulvQJBePT429ByoSXtLK5I3KpAXigXytx222QpA5WOsa+CDzbRRMJBSs+5AITmP923SyxzrQBkWG7WePsAOWAQuUuY5ZrbuJ+ynayfkIASY37XgIZMBm93KTBUL0abiMTbDrv6iPEdHB0xZXysIuch9GEt1XTM0xWrFk2BA2tMVTFqPgybLOR4ZySFUFMNa9FzxwIy1s9WwW/d7wxJ9IWvbNSqNmKkbnwG5uFsucsWpNeeaqcVVA1bjl7nP+woiGhmFARzaKRvg4ScFJbNv4XIQwLvvNLQFcx7HeHiwTD/UhsqOASH6nI4TO1gzuEvLxUItfb0HWNdP6KvgFwOhI8lGyJdCr/6SQAUhW/VnO9jHbWZNx07zDkWRqM1ZL5I9NudxManPIAmZn3Pixr3ZIvU6OoHp61gDR66V1zMj3bcvi5NzK16hJU9xP0G7EPQG19es05nekCgy3df5weWimZ0C5h7uPU2N6iEZL2rjA1R4xfVjzCf3uJTljnXy9VxC8H18NdhBKov06Eqm8eM+izr/pSppo6bCs4ajuXLpnldhWNuYmPwfSjlcAqXY+ZQet1LpANFV9NTUPpTEblrDrD6O+M4BqlgOSvkSicdZI0TmgYp93duuUkBVwizLPBZgZXAzLZTVv0o1ZUdtR+2sI4xGP/MBqTVbBoUanFH50uAJ7dg2zaIbUBR5sXUbN7EtUanXAmIbBqJv2prrsIFtpQhdc3PjSWCmz205wMzcuiApkAVJbdu7Foj3pkKTIIA2FApWGuM+lgyDdD1qExjMwyIxBT0LockCM42rwCdk/axGl+8hiUzKS3EXunPoN1mzQs2tCS4XHWXVcr4dARJRSFAjUo1NhzZjRgqN37z2Lhlnk5Zdrfhy+HRJfNF6It1BJH/MNZ4bv++TZ+hm7hQnsxyPt6ChJ8LlXqEKKtvmfURozlPTuhuGCE4WnYgsFjCAGpvfBiKVzbb/5FG6kyJFXE+eE7JuadFEJLwt/q6xF1+mfBkQXe/2pL8ihZA7fm4AACAASURBVAWB8iZZKL7apKtkrTk4HUWYBKpBkxnjtkH4mr5u79+oa9HmBkC+f1MkclZOpHuqnj7Hw2Bd3y3KazDj+rnK+sez8t+5xs5AVErMnNe3/7zNn88BNparl9mW0FrOKedI4aFC5HwNm7HUxqikV3Nt9b62jictaAiZ1fccq5OmoeC6updQ8JoU4DyRFqpa7EHMpMOQNdymXIN3h+Zu2RpumxIVe+T7Z43LttkqI51gqJb4PS3Y1xW5brPxRUONXjEZbOZElLC2Z7I7uUOH+SQPys1KGvNfJLrgvHr6FS1+po2EvE4Ns6dQAcc/JBuBMrbvbcqAfMR1MLYQaD+bit68BsBuwJxb1OWXErooIk4LTXgKaL88dasTCs+6psFxQ1VgEpHIckpQY3QyPPqb8G5qkYv5m7Cmzyq4jzDIPPhoWLgSbE4LEFVYjrcyN2EpsyqVjAEUAsqFcLSgFCPo3Isgt8OkqGJuCeUz2FXFYbPNJ2nMjuhpPThPojIV2zgtqjfrSyHdtT85BtM6cX1VOt7TaPkMHTvAd9EI5Hxq7wP3L9DfrutDOJtJZH9WINPRiTyyKlbZqsljAlz0136lVEZMmzIFSe4oJZHPUE+S3ZbvuiJAVghreh7Cb9wqkLEGIgLdTzq0LCKY0YMQ9Um6VryoIUx41txF1sv6GPU7jXIZ3T6XjtiobMOtHW28vKYCzIwnhpdJ1GXYSSP2LEaL7Ofbyy5tmnakEsmO26HhCzKRYDrxK7VlDIRWjcJWDFpVep5w3EPQEQpmLLtGeMDGLirZ2GcB1gS05av5/Azshf82JJhUaoNKUe7M0DN7pWdMh8FKWsQFWJbzmIBdl6hUuCmN9f/FrEn3MWBKo+WzN7UE9JX7voAYo1N5aU4OBm7pKsw1/PBy84aEKqpSZ73DOT8rRm4KUgyeLlkFk9Md01pYMWsqzpGKzTJ7Fc+fGLbLDF7LPI2l7iNPCf5TSed+CnZg84k4XH7IZZzGuozu+iZdW8tAFnxNoqIWGB3i0eQD2es1gvzO0oNFY+PeC+o7Q+6darQR7zPT1nABFY4BisdI0ac7axlQL6xg7T/EKB2Qm53GJuIdsTY++TF1Q/DCbrob69ol5O5xAapIJ1DDvvmgnsooAyL0Zy0ZJP1Dn83yd3+VDOguJujnfRQqcbRcbzG0vgdYpeieE5bVcsSZnNm+TNDRWul3IZqAegOOPQgIurBuoKgQ1qoFAt2YDXxtzJA+PAXThdYAdtYSYplH8WbraGmK1vwsfl2TOQGl7jyCg5EeTabPmpe57jUnzwB0WaY+7rWUU0PKomULErsEYdWhTs42BVJ2I2MEvClzWFSk+RkVuaSKQWIqqL6WWwAtusceFTRExc18s3iVtMYKZi0C8W4Lx4IPCllt3DuDakvoAjtq96w2gM0TSEUoBGUgyeMW6wc7KJ6BoRsAogQdAUl6cD9KP17TXe9PTaP7Yjg1xjoLhe+dqoHZDTNn0I7+uSC1WWwKArIoaMlUSgaDctXljFhkLYIJEouYpabNQfTKMFnr/CiDleDzxMQVN+HJ09Scm1SsuBBgwG2oj0MSBGk1z2uPzjXghrj8XApthDKy2uXpxtoJKgorAZClqfH0tLRnHl+HMxFGeyAI01kZOS/ttm07OrlWA7BcF7l7AMx43gW7o9NSZahqFFOXVBnUMGWlIt9oinQZFqENoHzrrYAxhQpB4rG01N1o9SThL27plTQzHWMA8UbQnztUymqGlkcJOwCi2SHUUPU4NEZblyPvOVHkhcyWsNlT8MNO3OgI/q1Vp/FYUpziWW6UFxrd4otkADCgyhqPOqZg0dsicGuQFpgZrPWZfJ+fWaZFO3I3KJhb6C53XadsBw9aIHEs2Lm79bM4gpb7ij5T0JKQssY+43jCmdZuqWvhXgvnWytQlX/ks1IGLug7JCjeF4oiSMtjlkI2YNqAxmXyIj6o+0YyzqLFFdEpKGJSMj70dwVgyWCEcXRLSnmqKAh24n5rY0rF1efI6LMY2ep3+tg8NUYFNxW4ZchCynqu0I7iZok9799sUZfFrWK4OhczoX4GV2NMFbzUHBj9p5WWIuTzasdsWHWXsjWZvg6h457ys03uG2MWG5dH6KP4YYMGFHC1ep+lQQwNVHGiHEN3i7mWzoOqvAUQ2XszZYmZizJS+Twxf77bOwRKzjRWRPPOMkag8sh1Ljmd8Jmfkv98IupOaBgnhweiuZCxLLgTulk2cgt37MyGR/+BWhyorVb5v462CN2XMlTElkJnLPXtIhnPHtTojHaPUZO2WiQJN0lMmOTcUIRgbo+sRtmdhkS0uF1AR0avGwFR2rb/WFo8WuWKhSX8l5A0l0YKJQvQNN68Nh6m8bG5r9AWhZrWR3QphaOYjGJFJdRjjGIUIN0D0qJ3ac9AnIXlkLVN4ncaG4WJLk6z4GR6KfbMhlXxFDMpU3CeCyzrCsDOC7Ch1kMWt3/ekJW27DdXuvMC6a5nCwdUSbbuaoo8DQU70NfrmxHYuA5ENa3U0LjOVnNgi4WmVMH4VeNkKpx+INdm/Y2Oa0q/R6+KuU4ZVTTZpLxoFhulSrer7c9CykrSYgd47V5lySh/euCqQfa4l1qrrGCcAtU3X9EatlgEexUArQbfyhJt/ND+/Jbf1zNLq1c35RNMkRK+6ecowdtWsAkSJ6qh4Mb0vBuW2ghGhnDCUlbBJcLKfSta/d4v0Vjww1sao/PZI5um0L81FIO2PTTVobn1zuiBRSwwFG1FNydtJqB+Ck258n+5x4d9G5piiEs7fVuWCIDiOryPgciMcalCMyYc694VPHqGKz53q3Wsk7QYT2vd0ZIWqlCmi+bxP+y3amPRWGOdrQ0hN6H51vSxgYwl0lKmxpaIs/QxpivL68TH6m7lYHxAx3O2oLR6Y6KMJmOGObBC7XOqyY7QFMfWUSu3V2zG5uHypexGIDt+30HlOaUYAGYfSt9uGTCZSx2ImEPPeIJ8bi4+o7WVPlVkv8x1Y06+D/V+d4wRBU6bPHCehQlADFhRc0JoEnTq/SRUNaJBy5ikgrAU7s0zOzzN+SQjKQWNFlCSlU8hotWVuA5UJK7NuReQ9XiMAyrFHRoJKpKe86QFapY/fu+CmAhP9oyC1JmK/JCIxdEguyQl1jR3YcZ7h4RlZAEc11I1Or1HhW2fxef32hulEPsn3BRG4nhVk7poFwZsW5iXxovGZPJ0ebrLXJP4rCqO1yJAKgta5UAIjd9brKGqZiHUqSwd/7YD6OR2dsX3WbtlUejTG19FCbeLL1gXYWMXBhlUs4z3cZxJSQO4JV1sglovvivykZj1QiDiECiNVy8L7YUWNNS/TqFqpcpSKrvU9hXXqFoJQqQYR/Ff+LOEgmWFfaPUONkoo00B1W7RloblhpuuLLrQJOLoNRpo5cSeO1GTelU/0GBdKJMWOxHTc1v4JhQG9zWFEKidqfQj9xK6jZWkEvTGzCAyqFSrCuicvvU2pkPGg7olcdq50mZldYF4p5E5AVUMbhod8R0zScoUZZVXK8h3ApFK4ciqklE9kQX7K9SaTyomoi26tzne+G2tmIfoNPmA/AzQyfC6dwFQ71TdBVsdaE4GphbdJzAdYwnlSAUhCfJaE/5H5ReZpFBIPVPD8RQvOxT8FDrNCmFuIPMwoLpvDJx3jowUXTMgfGYz3DH6UMa7sTtw80UaOKLrCSNTQ20bnrKT0q5exJ6LfUOMI4Jvk5qsdQinBaFf2JhVFtDI8FOCL0vTAU8iHGkZPjqfwdw/GZVFKAqK1Yuh2AyJ2OA4F68yGWTMRBWjgrFVMJUUkoWksKXP2mM06itqZJ3t+2YJklHBAFLOKnPvyCatN5CRbiIlvTcYj0GysRwoQAYbwLKL+OlmXiFwtizJSLTgVEjMaDUMQGNACC7aeynLfEZvikyB0KY/BTEJ5aE4SzyeLjKKH5LtB2tLOnSlshPf1DzjObm2TXQ0prxfLir5p7cHSD4ybRQMfiRPVj9ZDUjKPdY5Y4aUh+Shvk3BGoITD4ykOayCyUTNAyUPDG4rHjJkgyz7ds71KPlo8V3Aq+Y/x1M0W1oANhwxtEVX6o1BngLc1NjlApBpCuoJqqZFkYQ5ey0MPV9ujiEhXlr8TCWObuETaUT6JxuUpiCN3lgYlSqixh0WzYkJ1dhOrx9HgGyIkndm+qr2EpiN6ADNv1mDQJcl2FfMXIU5xRgg+EEwBM8dUWEZBcFXMLYTIHFNGCozmQy+pgFhxoXfV0TcfQUrFAO279s+HIAbmCo1W65SxGty3AjjIlkVel2EIkqhMgCZzM05t82ERffKWlCxA5Y7eg1YTGs+aYnNgOyibWMJl4ixKkFyQxSn0Yo3vtVPxD08Deqc2WKR2/8BsOJWfEuXBDXWCDoG3UdXFJI5KlZeH1XVFVRF6fmmDJUAMEP0tUhDPh3agiE0nsiv95xtzYJje/2uYiPxTNuJccH0YbNoujmYLhrgEBh4CyqmT7Ueg70lIV9eel8EVbxDxUS7aGRKi9s2NAk60U3YH8N2ra/GXDP8wPckvDIUpF/3ZXVa8HWDLHKhCN1inpb3zuiSzOYvc+Y2b0/dNkPg2RSW4/EJYMnrs9LSGYjMhWRKsuxjpcJIAzNts+7FNKFko04jbYsUkLJRGwtbdNScBceZhjZs0odsNMt4DwA1+93sfOTn5CcT/wQvTdhuSahckFw7R73WgYytYiQhEmx/slE0N3pVk+h8dj9mYBbi6kqQAT1rLQbhyCMcM34h1zcLqQaKtlq5pGuOIRAS4SWRXu02dmQVL7OD3sq802CGcqRhjbVw0cfFr1KccisYr+rL3quJexCZwfKU1xmb3NLiNt2Q5d7hH/NtuVBWgRQyrfRsbVmE/K9JEpRVj/VMN0Dxjx5YGYJXEezMz7w2nVHItWeDsJrpRKEVq/EO0+L2wF7l5pkatCaAQ89VV3ISVsgprSnLalUQlmNpaappoSji9dzxWDGTgpaFniAmgIQEg8K2bxvnCJOB2hbt9Rz+nRaszgzB+Uxi7T4GAa3FFBwAjqEGzor5NLgMyIrquQ2+03r3zVOygIB4oltK8aL4pA+3gnRVF2P6W0pmMHLDHhRp9RkM5lxGBabj/zN4yAD+bMpXMwqjMPK6qFZN193JJ3X9yGItxjvU3zZjMqzHkPyQJtjShGXm6mzFKxQH4vpQYTJD1z9fNdeq87EtL2iTZAZIfeVZpzuct88gYRkzD5Zni7Dc2ABoa/lcVauvc1MT6g4230jCRCASSgNRo/YeiGgNcs1JyCq+qTw8qympECDBrevS+k7616b76zmBGGphXM8XTAXpX3UTanQj2GnofjmhN0vnk5AYy0G07FPL9VKcm01yKQiDe19GBN3k/inNlmug8yCYNbA8v8JrLqAt3OWcBJARhzNPbBQxFb9cDFpMUp7KK43DzGdlX5Eaa/DGGEQtHCGaSzBKUNHWBji/a9bYZXUi3blElVT4UqqmOAJtbikBLz7U+4u+FEKxCA0KyohJsVFBIPhCsZkZRWrdPemdv3scgkw2xoEMWCHxnnFptROikaly08W7I+26IYKUTXGfCCbT7fN2nkwgYja9WnxnQO5sCasrRtF+/ZbjZlAJqdnUUj8nlP0mVRadPnBB8OaKbPr8LYDvpagIm/RDjZnPjCROwrIMmpIxO/PHGqZF4J4FBce2kI+t0GKajLLHFZ5NWZEL3wtbtF3ZmnUUvRzux1KwjI2oQc7mLIuZU624hMN1sFOvqXCdVD8zwzWzxVoJhQ4r6rC2CFq0UWu3Wl+NnwqUFskAnfbGtnOEEFTuVLRJlzg6Md0Yjj93n256S5plGhvp5ZSbOMYOcz0upeDMPlQFJ3LOELJImM6U5QieMmdsLuc9t8pJtLO+zi0dm/tdWAchZTrTHRKymqg2h8imP4aZcUHxLVoqlGuxHkPZn5yPgVMa8HlUrjD5BVkzQrd5GBzMosR7I4BdBXvItg6eCIKGL/ZGMQuVaHBO28Esznpq1kOMIo3PirPWMo8EduaUd2KMSgsumAnZqbV5b9UOkBFZC08BbzULtHY2lBUglOcJTeUJhsKRxQZSKxf0B5vOkNmaGBnPeKXgB7tC+zKaRVMl6kgrLfg4oS7PMLCZyBDiSYvQTomqtmwVne8ZFIxs4EJU5iVkcQXTcAXfq1Q+rB6rKVhly2vp28d6F/JiGq+XwNfGtlEWVBQ00Upo0hIo5+/us/qaDBeDEv1UGq+QAdD3lHhYZqI6WPEOLSw8e0mQD9pu2GxcwywTe6tCSt40nghMZzBTNQyLaNXjTZEuDZcmapTYUHcVXxEleiovuspA7t3gXDCgMgMUouGaGSzPbwWMJ5QBjbdC2fesWV6QJCKdaDAz4GxABXirXUHWjPhOVntQUZDhlpxovtg9LCvdgo4OpJnoH2ewCUirV+dWxuMZRCGLNa0OYEix0G9u/n5OWmc98h1pJZXWdFrGvC+VnyBkLBEUxEpFY6APiWJWz+eo6CgWLNzw2foaeCglbnzKQKpYOBVcWagedG3+vJBUwu0MJntW+JGucf2yvT9T1BUEJQJYReeKQ6USSqQRdJyojt30Z5lrb0Vpvobi7nEdS1rMrLDUuw2BHPkuojvX87n+wX1U7GRwuhUu9CIEZJaxnFKaMmDWU5lEWOzmbVBFalN3MEA1JG39Og/SZWMhl7arZxwmmuVCBi2UIHdz8nkFlMDYUAayo4aj0Cp/V6yEsjeWRutcCzb7wdjQd2z4CqXME93pgOiOMj3roYZFNqQCbawQawSmVQBkBcsvrLZrQfy0vNmJuqy4tYmS0TwFFah8cRGu/Cxa2AXqlMx3joyzsAGKb3e6tuVH9SDMvDUVAK2tM9/PRWtWBJCVCyaMeVf6sMcryG20b4i+DPMorR/SiiNoNSAYysyRcugUMjIbT3tTM5JEDowftViNLIdR7bXnJPphmo/Ww2lNnPzAeIWh4Hjvv0Drw/HSQud1qqrs6Ky1rKM/v0lxlNIWn7i3a0zz1HPd5VeHAobSgKpnyO3/jolBFzb5sfawROCaGYrUGnld7QAFd8f6HoylsX1A0bhzX/GFirm6NIjurk/VByN5xdVEms9J5AIrg4nkpbG0bFohV9d6Ja82pFgNnGKd+tpKN9jwXQhW23JuPWhnGyEsOBSLNLRjcUmYxgAPFQZOLAh3kw4NFspMNCvBCYGw08EOyCJ+i9jr+Wz/X7wAlfzSYvoaenYg96YwGDvyvlbtmNoe+f7ei0LjriWsIwHHIqVUwptiKzhbaErW0yBLVL4/6TXB+gnHVklU0dSJTJOYyzb0jHG0TUwAZATUfoBCZsUX8HJZsk5kGI9eYPCOBXyM0eS7MqoOBYsrXtKNEMvKgxcoDC2r1WJSxGkdcXY0Udk8TnECS1pXxh2kdKb+ll+vGEQ2Qx7k06ng9MmNWVLCs+1lspolFWL8TYFcar37xVy3lpk0o0IdCm6XYV40fxkUawKPMF7JACCTS+k4U/CMm6HdN7JTVg54MnrtDW4yuGOWTVMgAeqblqIxzoqxHIIbedSwJaFQdKNu5axCAMksFEQn04VymmrQggyYEjZn9DbrNXw9Euxi49t4dLpJagzSMg6tg3FEyPfotRhx5slxODdZ2KTglpRBS8XZAl9XPYMbyZwLREtJhQM+Zy1hTHoUaqlipu0GqQl4+atMXNfzUtn3GA7XOenvUm4VuAtBzI7vG3eG9QKpCKZXFXHji4l9KpF4dnTlymd5rk1CXW8CHsjDxczKpmyuq/hKBU0tW95tGwMVpVLAfeZethXcSs6dwW6l7JCxh3hOry/ZSwk4i9PoRpDmc0bNMY0jFcR6FNUwPjGZqk9U3U+BIzKpZlTJ836yUNE3hhwI4zc8kNOmZL4dAM1OaX2TGpVLrxoNOaDbYpjhhgTJCMUJ/Ri8StdfRUGybJsfx1hORWloEidQW5SPVguzsJqebc4ANqcBasceLUhBZMCxZGAo9tcwjTSCQGNR5+3twUIkPsKNskz8WG5uCo0TVZ4MrhowZiEHy+BZnE2SaGFC49fmMSEQE6OL6d1lsXu2I8bVlBqZ1QC2Y6uAVebvpVz4zKEFPd/SAaoI1FLNrHjkei5V/2AjPd2qKeC79fsGCVKZhXAMG5g+sVgc0DTnsRoAc1uA7utZMgPm9ArypfZxuppSsgB96zF2IXScx9hJ4CnkGrMDLF5DupE2lnYM5ahWeKmESnh4KFW8MxRvvEv7ZgxAujpYlpxn1XQAHq35xhKfIwO0YKZji/xiHTNQ7h61No021Y1eKgbqNnYeH1ZWxRKlFC94pcqtnhHPOUCm2hJpwHdzrnCsseAUBp/q/+jpWHkyjSrKqEXy9xXnwA7bRiJYoILaHFVpHMKbte0ErDgAo8SVVpzGs01Yy47S/tzklSd/QcIwAv62vLcY0evMB1cgrogYxV1pbRjvyKBq5b6trBDH6wbDqhSZBHh60jKP9wODnITiAFPDRE2goIDIgTJuQhIddgtZoOav1m1iyGQSWmAtcjgdpeS6wFFpIy120Dt2AVevhbmPeMT049jCP/fwdEFCI+xBBVsb9spnnOtxCnbFb1zXd/cUmOtxfE93BaRvWtPsKan5qZ7ANoisrO9J5Eb+n2DlpGM0HmClL3mUyiwzLIlMgbh3rscYfJdHSrkQ9ZJBVSTPZwtAUmiuLXNXSNRXup/AxAoeu9kRYd8bVeOkgqFxsaQLCkmt+fdMwOCr7ZZlB/cD9EKZ2uDCRWDkHaHxjHB1W2Pvo6L3ZGRI+xlY/jpyo1GlN7O0h9A1sw4jNwnN9bg2d2FgjINccN7NQ2/TylKzpiukgh5vY2m/8+/6Sassnz4Ykoowvqcg5zjaQnJUAKpOAgNV/htMN9K37wKudBdjacbmQPShm/uCeu9mrw4QKdgs0KlAbSkLvden6hoCbTVFm8xV8JduW8Wg1L8kJlsUNFMjYirreHW4OUSM21hWxktQgVlaZ0H0ZOZqEL3UmlDwlD2oDJoyVuQjWnSiJb2v6hp61szgQVNSXugSUr4K+nsbe39GrpX2rQDoMbIew6lqUJ4dO068j0Hdip1E1TU3dLYAt5DIrlDjJrCcNEH1Eh1ZlBnTHFjmAXY+PWyKJ2roAUMSMK1ghcMqwIJ0W9B+ry2xgPWJKlZQu0Ar0FKpwKgYqykMleOiFpKT7Z3JFRAaupfPFQPzsFyVf3P8JgOvudO9yBOkuNgboQttWIxHd20sssY110BMwxbM1n+S/NWDWNoJqbkQfQSDkQk0To0n5zl6AI8WzSUEhKxlSVNxbOIEBctjBFOKSUakuQmR4ZgJjwfcjwWftenMSog4IdWVAMVHSVOTQk3lkhkZrsNm/vyR8JqEcdM+UAos0SXX31hXksG9pJwUY64CYxWb3bG6ugW+abVtQDtCNbY25qzyDdrm3FXTxPt3ol+nPQPNJ89qrZghx9mRRfGKtzH2lHop95kb8yZ2rA1XBSThthnQirDYVwApcAwGUks7A0fwhFioa3r/C3dM9mogkTbM7hEgJBOcDOyUzRH8LoXg9R702IoXUyjQdwKyO5mC1oYoZdQCtPfnIDJynjBA9yCFDW0RqIxyqx0XpI1Hm5wssylURHZC8BXcCmtUOyCtDUyaD05GAhVp0plm0BVKi39Zhs73SniBrijI/D04zGWUUK1F8/iOxUpBCWfdSCqdjb1Ll6f6dJBHjBABAcK8hBolqDVvJJzOuhZ4IY2O7JowxqtokdN1YTxgmOa4Ha6DQe7ikXQZFUBuiYHNzdwEl4qWAcbGz/quBZvjM75jwhyYKORVcsBFYSA8eKcHOUFl5VU7xCzRAsMOiGDLeQcQgyihWYQU0JHVY9RkkRkYUaRjlb6JZ+9K06Z1tVlBQVpkBU5pESi4qpGgUA0RBrRINjCxipxcYBkvmAKpUihtK7CZab9GWLOTsJpWrFw1PQoAqwkVjTdE0YwRHpuYUqFDpiaJXkA+PWmtSwEo188ZZGDvfMbP60dzEZpljHVsFtCKITdWzydOVu1uxxNiqoBpezdy7TYWtP8EPNwE7gqG5xg3FnijzqC4hzsmN0NZ7R+Kayr2JetvnScTJTlQBweh1iRjU4qD2QCMNQmjjaoZHgUWWU/hffjJR4vSnoWId5tnDDuoLKDxvs7bvqHt5myVucqA9WwJz+/pIYdQkmwpYJge8qwAb9b1THfsLJlCN1v/O2sTAKg+wVBVhADYbaigZSABCY5PVFEJNTghbkYBuJC5cLQ0TCP2lFgcHMyNPoaZe/dr6p4AhntbyiKWn0iFVMzN3XVSmCKyw/SuCWvvSjMFuV9cUC8Ljex67gp45lucrO/JD1Z04yaeZuV4U5Vwm47HUxyhXWtAHlZdCl8WXH50Wh4pg0SP2nNh4JkREh4+PRGj8BYFKguJBmtecpZFa4f7SD1fBV+eex3KczvBJ7SyuSY8WDna8te83PfKyhShJ9g8J9h7BRaaFsuCwxM1J15xDBkYr7oTV7C2lbxbpNktaT0UzwuBhNdxG77W/hNv3c9ZMBj8U/QjPTeyAvL1UsYqx0m1ynV2dx303DzzogE8UXIiFsvOYEk/g/tOPKOJ50ibbxkTHiUcgmbJbI5iJuPL6wyLfpR7/G8qHYqhnlt/c5MQchFqLOVjAQyWDlQ5bU2+GzoSloKNUazRaVAMxnnW9l4DBCV5HZVD98NJr4gFARspKFlPhuyWGpjW3BqYGKqjh0Jhy/b5G7RHZq20KLj4J+IF7sWkGh+aFQfHyToHYFOhqfvDunu6WDreUmubNGW6GDn2/Lp8//a/RF3t/virI8Py1ylIxnXk9+etFSo+oVPYeH8jRPM35Oo1+sHRts03K853cRqkhVwjxqI4diL7kUOgu1NrP1rFMXI9hAQ3McaME3Ee1mXMG+1ofGqtJP+SIZdM73xOY0Rcpbue25CtSqy1taZ9NgAAIABJREFUc3ITNDkhXJ47Igd7bgbB5nosaBdpxFU5cW6O8ma9GJyhFffpcGvBKVpDPs+j32HzmFKft7QW7zs5ZqRr1Y6Dc4SlG9n+nb7unGuej5LjsNTsLHVuhOXeB3c2im0dp5yIzcFNUYTDha7SQmRco5/f4WAAyrLMgqXNwXhUpERYQfstqtMaoqwJ4yYGC79XwbRWEMV4ifdahJGGrmIZ5llMx6AwUQyfwdgYsHlHKSmilMw4BbMk+dacNw1RmcpeKBiCmkLLAKe7lIPpHTlCIWoqamYTshqzZeu83yd+arym+Efxmom3p1KVm/viItT5HZ4CXTTT+BKJ0TTFZxF7qIJGaNwxjFQMrQWkdv72OAs8vQfP4D4wfW+7MRZ37CraCkc02EUSI63kyUg9BaJ9Hs2rYnddt8C9RdoYuyxuai5BfJPvZmwCutfSStlguzQoas6U1epHqfkrEu6+YqgsNjRw9BRkzKRkt6xalhyPbRTazIIxxYS5EzV9QLW+Y9AyDzNSL4rmcvm0pO0Wfjqfa4SrI0+SqjSkmD+tjPoXILMGUhrW1qsYYduujkI0EwEeliWW28GFyPGynWEy2RiHepcUZd7FXiZyj3yCvVPCGOxIfESWiNaW35MXOMcUlRHIphfoSSDzmVPWeKiRE6z6Pdg4iE7xiWiCZygCLTU7RjQGtgUsqop5V+2HwTalBqPHeVLhmkXKf2agU2vElvutFqKjqACgBsYUSAU37onyRmP2ldn4cyjXdwKZclXqeLfb8BWSP8cSR37OpOmYB9idjKwCALt0V3CntG4FkE5kIFDauVtwozTWX4Jo1Mw1oUpFVYViinAW06g2gwHDfDar/xiENSwFt8SA1LgTAal7ALHG1wncO2YDFTSsTlKFKDQuLk7SptJmU9awfHC0hSyG47Mi6NYFt9EH/aesWLkeJ9AFv0+ryL09hRhafKKVG5OusZRcyylFWtbc6t3jAO6tL0PNFIzX1Oc1505/uUdUQZ3JeT/dlxOxAx4SXPtEOA+JYI3Kvb23ltOJHOnmbAKnTeC9ZVq8riv4z/GyxoFHaNR4NzKEJi+JNDqf8n3hOVGmtqzQ4zwbejcF19HsWA4S0JAf6tiM/MyjUxb7OxjAXae1WKgJWxdYKg+D2pbl2Q/suBQTKyvai0eobTdpU7OASOzpQOvS256B++1zSKKBY1l2GV/rC4caKxgENC26GMWRC1NjAVzPt7x+2MDKbmGyWmzb1pTMqC3F/X2l7Iq+9T1L4a3Rlj+8jyhhFg0HmwFBtCp30duz6N5VvCFK5R0YVfKMtJQFzdOSz32eeJZj1jsIz2N+k0V9E2B/EzJ5wWOOpwzENnPim+dKH/csknhhq+Qnaz1OnJEql9onBmrXtBYYVu6Yn3AzeCVjHpSVpPtIZBH/DBhaIymrs0d7GrziSNs5sNdrvTtrfIg+19bNPflmzlWfbRWtKK3fKquWvDG4WWyJ7phwZVeC7QwDI7MhYBTcUBHXwgHlV0FCVD43Sdksfvrp9LUD+rUTwMk0QhFZS0EI2C28U+gp1C4NYY6A+Dz3kT4+idz9PPp+ZBhADCP047Tm0PvYK4A1Aay+izhE3euiE/3qKTdBwNzDanSYWVofGqPOuWyQlMhI9kcxHm/WnsLQNnvJFw7tKswjFxLbH6Itd92/OQg7laljarNYPN6gzBfCQnFHKgVqW8zEDuO+WW/RIQ3DFpJzTonCpEHKAKhc3U0xih6ohWJXU4oh1iYVapt7VIC2tWFR2lw3iMlyvUUf1SZxKwOSX2wzjlyJsvL5w6u4K9rEG7LeINJ0n1UF0FAlxxxM3bfc5xusyhUC7bYwhO4lP8SvUm1VmOHhy7VAFmShS6Cr4pKLlYvIAI+N1MKJRmSNoGs6hCVBKDAk3mRTHX43edgL7/NSQN0OcBxOwGO1SO09GwKB7942KiFcFEuz7R4oIGt9R0FMZSbFSSvchZPjA4ox+5hmU36NBlp0pjV9TR3u7fo6EQ3aZVmWVUHi3q5v1ruiQTBpzn051QG706XG3GjU5mJpUc2KX7hmZYg8xsJNbQ69n4HeaNOYLd/yczVo4d8q/66xDY2RaAwa0+b5VC7kV/LITARDepIbZHy6kJ0ouNrwGWlb1zBjIT5Nrq7/LSPHcVkq3s6nnEPRhWuQigolP8UnrkyO+wzl1GmL0gGBxjIoYSJBC7zZyP0LkoPNzwZ5kFZNq0JW4+QDHITRm88NYMBzw1QnX+wNtvWUZdfODEA2a8FhRLCJgZ5kckF/umUcBNNdaNe1KYHpW2DsTuMBX3UVDhdC5fMtZhKpPaIUMRJ6S4joovjU6ySOm2cAmxPellN4xtO/CVecLtoyfiLmKkLqc7PmOLXYCxEXIe7Fl12Br7zX5yd6aS4jDJdccQXue8+7AABO3e4y/MB3X4OBtRRcC7aVC1prV9WStVbwgMiDropxPn0pNuq83kfOZlu9jhZyPJat8ETjNteT7lEPNBI1FPqDkEDRkvd7G+GW773Nt3ihre6sta51RBtXV1jdE2BhIwQGmAGT4W480ZFVI5BGPRAF3qBgcoIQtN+XFuJ1RBeJMIIwDBiFRuJZDyxeQesRKbgWlCoG7YvcNCaLReoczbIkpd1RiwNAuwxB7Y0iCN/jcdALFeSw2DBkFj7aSMaQMNB65/yogWk5vvwhD8KLnv8cPOieV5TlzjFo4dpYC9X0YFsxRqdH9SegdUy4rFhBLarZDg+4/71x0WE1LrFkOq1vW9P6zGt+ijMh6Z1Wa674gqu+DD/+vdeiECPpPXH3+90XP/rPHgmD4+DUBXjw/a+KbVjeLNosq2+kOYWBe3AkNDHmq776arzi+c+IzNiG/8grmQLMdoUygEK2ndaW61fzpiCNTPWGjFX5+UhFQ16vtaIVhtZDY2ryw7nxx7zqPgZRVpOv+N6r9F7IlGvUkNLGYDceVzghaMHjCOJ9a/ESmsFIfcP5cK4hE3mhNG9qbp6iFRY4oV0LVPKIuvOPqsu/bbu7lMEexSpGKyghX/RfNF9r2QMKA4OH7c1dm4pVQmt7Lmz5p0WAvnkmPmcgqbtgLWPk6ctKQ0P0+NbHPwQv+rXX4omPf2hTTKWlKdiDBTijMWCzYiaLr1VTGrJbx8qyFKw2AFjP4Hue9VO4/uasCeAY2fSXCC7bFcZ3hSAt2+KVwmAA27JepK0PT7uS1WeExnDLTTfgW5/1X7B6dmgietEmOyK+ulcl3ySdY4siOtKUYPeg6ba2Rs8yQBXBqttoytsMLmGvhk2b7d2gSwZok1eOI8a53ZtC2nUeQN7FXrFCJ0QyKTsQPU5k/9LYjpTXoQ16tatVMiqabWWwZLJtu5Ds55ib8RnJJ7sYIGsWYjg8twCE4Qa1fKugW1lrLtzGn3ZESy/BIS5yBjVnixZz4SjEaGXA/+BnbfejtwXK50RhCkrD8jnuTTkAaNvtubXZQJ8yFkA7ExvUY3Uig6HuE1d8wRfhXpfcgm/9r7+DF//yc/D5l78cf/vJ28CNP9/ybdfij1/9Ohzc8S543Nd9FZb9WbzsZa/FR/7+Flx5jy/CtY+6GofrOfzGb7wKH77xFoSCGLjv1ffDQ7/6njg9Jt725j/BG/7kb+AwPPDhX4NHXP1FqLRbpAvf8JrX4Q/fcxOe9t2Pxm/+ym/jE2d2eNp3X4OXvuh3cecvvgce9fD74oJlj1f81mvxges/E+SfwB3v+nl4/GO/BpdfNPD2P3onXv/2j+Lp3/VIvPiXfgdn1ow98F3Gf7hmdNU6SjJccPEVeNa3Xo2f+cVX4/B2l+PJ194HL/7Nt+JRX/9Q3Oced8L1H/owrvudt+Azt54Dj3i415ffC1/70C/DhQcD733Xe/CaN7wXl155dzzjSQ/D5155B/zYc56CN732DXjDOz4CmOE+V98HX/vgL8Myj/CmP3gb3vbuvw1VYIYnfNu1eOerX4NTd70bHvWAu+O/vvDluG3NuISVzx8BayoP8rRLYfDUO3LTFIpJfpyrjOvkAUJUMR3Sb9zknfis78hNCAK28adoVACehizKA5gZivLxjihKCcavVJAyuWDAVB5D63NrQOuwFp8NnxXYmpljnetxm98aNeVS0h3yAAX1+Xs5A+bWrmv/JXN1RSBI7SXgpaXRPoOuSeehkIaenzEJMXHzWZMAI8vRY7RD/8fnAbymdaxyzq3FMPIZj/uGf4JXv+L1OHPLZ/C7b/4IvuER92mWe8FDHv4AfOPjH41/+bRH4voPXY/b3flK/Lef/3488KFfg+c84xp87MPX48I7X4kX/uz34cLFgOn4tqc9GY9/yD3wx29+J17/1g/gyd/73Xj2E78aAPCB934AL3vFG/Gyl78BL3v5G/GqN7wXD3rQffCZT34WjoFrH/cwXHpqAOMAj33Mg/FPv/Nb8CNPeyRuvP4G+EV3xAv/yw/E9w5cdb/74aW/+C9xiZ3Dn777w3jQo67Bjz79Glz7mAdg53tZZMzY01DZl1yR5uZRecAdhxfcDk983AMxAJy68FJ807UPxU/+1Pfjqjuewp+++4P44q+8P176gh/GXS6/EHDg/v/k4fi3z/w6vOOt78KrX/+nuMuXfDn++VMfjs/eeCPe9CcfwM03/T1e+aq34AMf+SRgA8/6oe/BDz75IXjX29+NP3rnh/DEpz8FP/bPromNbQ489OEPwBOfdC1++Lsegb/98A04Xq14huvfEbIj+5YMbJF28MXIw8A7X4kLGm/wP3cPnvL+3jSqPXsi/gLYFd685CzISmWNdJ+yYY7Hu3nEQARkPZ9DNMXMDuoz59rNJpsxrgg0I5TkrKrTQBbpI7EoyDaZjoRFvYw271GhqccMBl2YTNsFWCAsstSMsYMNVmTvAbJCM6wXmPDcUUpLXtWWlYoDuBeiEAfVTa87oJtRzwDMvP3NcVaKd9jAMMvO2gzqDa4yDi68HI958JX4wWe8GGaG//WKN+CX//1j8YLf+hMcu6UfuMNXXXUpnvGc5+NoBX779/4MV7/i/8XTrvkiPPtHfgFn9xOvePW78BXX/SS+9MrL8Y4Pfga//sKXYF2lAfH+j96M//m878CLr/sTfOrjN+GTH/9EuCfLgh//T/8UL/qZF+LPPvRJLKcuF1PBgdMXX467X3oW3/Mvnod1Av6KN+N+1/0c7ne32+MP3n8z/u2/eSqe9x9/Dte96UNY1yO86vfegm/+zifj2gMGBakEIHrc+aqr8DM/9WzRIKyh4/I73Qn45F9LKce6xHPu+kVfiP/43H+NP3rfjXA4XvWat+J7fvhZ+JFnfj2+7z/8Bh7z6Afhpb/8a3jzH38YgOOd73gfdrsFcwLv/+CNOPPZO+NP3/VXcDju+7B/jEdedYinfO/zcXYfY3vrW9+Ln3n+j+Efv+U9eN2ffhSwBf/oTgue+QM/h+MZtQdVB+E4GZOoyJGLZ3plaZyFk7+zHsY9S5C6i5wInYHN5mYSlpG3hxoDneiVkuOgPG6aG2fMge8xG8CMDXS9PeDcHKDE2bG+Kf2Dyac2JII2bklFblEntAabpioaT+HIAFDbHi0vhO4J4f0EMDIXnf52/J5uwDwG93VQOWz2NjgArHIBYpGqHDYCihmYI0RqwcPqxLRo3HCW8qaCceoJFymqdBdqLLstEtoingiIhf/+FQ++P25637vx8dsch4cHuPmGD+ODR1fgofe+I37/PR8XtHv5y16LozWEa3/2Fnz4xk/j9b/7BpzdR3xkf/ZmfOijt+IOl14E909i3U9ceY+74Uu/+C7w4yP8zQc/Ab/4drjg0HHz2Wz15iu+/VlPxdm/eBt+43V/Dri3BsfZ2u7oLF70K6/CPhGi+8SHPvr3uOIOp3H7/R1w13ETXvmm98P9IJX/xMuveyN+6AlfGs9IF4GM7AA+/Xd/h1/5768u+JwG4Kqrr8bj7rUDs2EAsrXiirN/91G89X0fy23QwRe/+qLr8Opf/V5c8JO/gfe894P49md8M44vfA3e9s4P4KZP34p1T14oaGpmeMQjvxqvfdXvYTXDwYGpTuC6330Hvv6RX4HXv+tjAID/9YrX43gaWBtTGbMS6ljP5u6iUvdxXxxZoEBjz0Iwe+MA91IpeBnMm2w743hJKd7KIpGvxWNWdSB0KXhwc8lj7eNiqYMjWxPC1SPUEeXlHCfrR9joqg5ebhWlztIIk/zC99oE0oKISUqenIQTCEAk5sK1rb8ZdOPeil6KLV/IhrpEqWS5BVdYzAWUS8MINeCYnv0TUmGwco2QjczOhRgZrNnGNrzFTEKhUCO7FtCb5m++eP4+mqZ/0jc/HHe9dMWLX3BPqZ8LLjnEtz7xkXj9e16SXZ2Bs7edgyAhgON14szZc4CzwGnFejyzT8UBfvjfPBt3mDfhla97N44x8MCHXY2LdwPL2MEssg8PfvQ1eOhdVzzzR16X67jbxIKipNtx7hwbDsWK7teY2yWXXIgzn/0MjqaBBwmXy4WkfxkNSzE7c/PNYeVVA5DW8nO+AI/7kru0mgF2OrOAzbaAoTrAce6Wz+LM6Utw4TLwWy96Cf7yXffG1z78fvi2pz4BdvZm/MLzfh1vetf1sm7cfn77yy7EI570TfjKR3ydBIyK68/f/nYpquOjYyjDlMHlKHZqNgOO2uYPCaUUAuh2kw9cAg2Dji8YZtqTIlKPge5CSDnQ2iZK5z0Q3QwVj4rrlDCAxxYVrk12kO9xJRUXdp7XWpZSgrc+nDKaaWznHiylt5kVnIwEcyv5tBJsLkLBm1IYnPzGAjuyu3GrjjPDQPQG7Od6EA2oIaueD7m+xYg1damr8zIOBdk3/Q+Y3mzEGMPqe1mWtHiyPhM+Gbit6soIloZS+5x/dE981Z33+MZv+Xf49NmqnDy89I545f/4EXzBFS/Hhz9xq7ihxmtSPhVEKvRyl3t8Cb7mC4BvfvpLonWsO/7wLR/AU5/yQFm5z7/nvfF/Pul++P7v+2kcz5p7uUijGIMj2Lhkhr/7m4/hgs/9Qtzl8lP42Gc4LsPFl12EYTxta5UbWXTm81iS3T7PjEfNORDjwcW3w8Wndvj0uRldDH3iTlfeDac/+b9xc7oS73vXn+Mv/uwvYAO451dejZ//d9+Nx33Lc4u9ci3e/1c34Oy734//8ItvPG9+sxc95Xh9wyM8I4TdzPoTStipILbNhePLniKdMpYVy4n+HKMUQT5bq99kxhMt+ebacgk8mzJB16V7xI12UixIJXX+NWzjsFWClnO3jXxPBV5rv42NxQfc3dx0DIArF5//McOR7eMqKBj/1fEBpflZeajqRAeqXiJ2VNrm/8ovQkK42lkxsiCnUkXWrB2DSyO/G1gUY2BaadgOY+yEUOL7XTxbfw9ZnmELFlvCgvNdGgevjd8f/81fiz981Ztw87ka9cDA8aduxKveegO+6evue6JeA1CgC5X75rgsF3t/dISLLrs9Lj69Uz3Awx71UFxqceeFl90B//e/fhL+n594IW78zFEF5kRRbOCwPvcqDjI4jj99I37t1X+Nf/9j347PufgUBoBLLr8CP/jMawMB5Lo7j2nsEX1UAV2w9Tj/fYDqO8apy/BDz74WFx0EGr3wksvwo//iSXj5b74Oqy/4umseiItP5+a01XHD9R8PMOwGn8AFF98OFx4e4HYX3Q6/e93v44GPeTTuc+UVWpvL7vh5+JmffjauuPCwxqZ17vU0B8VHsOSZRbUUw/J6iyuW5B3xjHVeWBQrYBCTPDLEDxU7s7HoeSUzO8AbH5IXkIjYWv1T6iwFWX0rOyOvqWchr8szZrP6WKvj9T1llegRDgVn4bE33SILsUUHLs0WD2Mqh7sjlb6kD2aMU2RnYAcwDHNd04ozoLKmtqQ/BsgPdLonE4o29xSqCqAABnlqzPTVY8TbXZn0E8MS6nNnN2PIknA+LkQ1Cra2lJoZcHjR7fGEa+6F5zz1vwGyPgyGTVz3W6/D8370GvzCS/+oiOqeCCsREKbGyq8B4MYPfgD//Q0fwYt/6V/hHe/+CC67/aX4yz/+Y7z+L8/iIV91N9zx/o/BlVdcgO989lPwnc0k/fav/xZe8/abig5tI1WZUddw3Vf80n9+IexZ/wd+7SU/jps+8Sl89tOfxvNf/Fo88t5PEJ3Yj6Nnq8q6xjwEmx0ZH+jWGDj3ievxynf8PV7wgn+Fz372DO5+j8/H237v9/Fzv/aHAAyX3eku+KVfejQ+8jcfw2174Eu/5PPxsz/9K7hl7/jIX/wNPn7wJLzyt/8TbvjrD+A7vu8X8EPPfSn+r5/45/jE9Tfg1v2Cu195e/zy816KT952DMa2at413uCvbJoUUlxzoEAyeLlRjhDPVr/NNLIMQnp/Rt7FLFHu9nWemcLngKi3ZKnkoO1qbXzLsUVsA8VPGjPRTyAK+BZd1fMo7BUjjHt5ZcqiO+ye937czY4LL2YAkdCj/26dQBKIra9vxoN+mKqsIpeKDXSc5bruJDTetA8DsDmdbD3GsjvVngF9ruPc2r0ANocczeyNOHjSN1A79sB1XWvR0seNQ232Bes9iqouOL3DmTPHjdicT/x+4YWncea223Dq9IU4PjqH/brPwKjj1KlDrPtj7Neiy+HhDnO/4jjz5rf/nCtwxaUX4IYb/h633naEg1OHYanHwG5nUI4++fLo3BGO9xMXXHAK586ewzonLrzoQpw7cy6zUMG8p06fwtzvsV8ndsvA8X6P0xdchIE9zp07xqV3+1L8j5/6Rjz2iT+Bs7PclyiqGjh9sOC2s2drvtksZXdwiMPFcPYogokXnN7h7LkVl3zuF+KVL/gOPOwbnovl1AW4612uwM033YSPf+pWwA0zeeng8BB3/rw74PQCfPT6/40z56ph9MHhIQ4PBs6eOYuZG8V2B4f4vLveGQc4xsf+7iYcHXMvw4rTpy/AenyctAxBZq/VMXZY1yOtJ1vf12bDxsNZc7TdBVtuKRTfioOVavcuQLniprDO/z2W0V3qoOeUsNZz6LKv7d3IeBCPSDhRoNbaE1S1L+WtXHiT0uNcsp/FPA5+9Ztv2cGnTd9jWFWH1XFm+/QBvQSBAp0vmfO4jmNDuSNTmm4FW+zFoBDH2SkbUspJ9xsnRiXDoAsVROumRbrougkgOziBkW1uC67sCRk0XhvaM+bBU804W4P2sWS2aE5WdDpuvW3f/Hn6lBV1v+22M5hzxdmzZ5r2DwR05sytWkj+2z/z6bjp4x/HTR+nNTQcnTtbCx8cXFajOeC33noEWrVbb/msaI1k/jO3ZUfwscNzf+r7cd0LfxXv+IsbsV/3OH3Rxfi+Zz4Or33lH+DM/rj52Gn9puOWowoCOoXMDPujszjyVT0jbzuzh6ycRwXkuTO34q//6lbxB9PU8Injo3P42w9f35g7rZoB++NzOD5CGSlM7PfH+OhHrscmep+8cfbsWQkD4xTubPjMHpNURj3jAsU+bGME0trbLmUjeUOIs7J3WgufSR9uffdEakubf+dPaAx9455bZT+qFV7xt2StHXVR9DAZlMhejoaQsuCunZjXFeKcoRuANUwcuzP3CH+gs0UC2U+F6jHF8NHohkxE2nMpyCbojYSGOYE8rbqgVhLAdtKSYP0DU0YN9irtZFROM4NxhtpD4o0RvS1sCnaO0T0UGBc/RxjR+8Fc/NS46f7UmAZ0WG62a3OU20T3i8Gj2rQWV4a7sOpva4JCfMQAWOEla5/nXEZYpMjgxPPDENAqVdUe7zU4fvZnfxM/+pzvwg9dcgrnjva44PQh3vq6N+LnfvmN4oXRLKA6gRGKMaJPPordIKLhGDUPrUP+bggF4uD6lMBzngqKN4Gljw2d/5J0GAwI1r4GKjIaFb5nu3nNxdfeUozIjIfWBKh3b+A+5GKMZWTQc0T7PrrQrY0glSOFebvnhORZxWPlyHe+q4xhKBSIPtU+IL9vQhuJC4imlCEA0RlsLSPMz4cNty+592NvXufpi5U6TQZg9VpZw2b9aW37y1ITD97XFupkfXz3qZbloE3Ki1AU9LSYluPz/6+ut9vVLTuuw0bNtfbp/+aPRNISRFoWTVkKJVlJDCNBgFgGDCO+yEVuDOQmT5AX8IP4AQz43gaMXAV2gMAxYMcJHDgRFEWO5diSLLXYbLLJJnvvb83KRdUYo9YmvRunzz7fz1pzzVmzatSon9lWS9aUm20gEU9QLyzbt1HY4c5argFwmGp3/j/rV3hE3+xhYPTVfSDb59VRfns0LBkWa/az1EYf8LRgHyMJ2U1a8er50M9vF+vWYWy6j8P/nihk+t/IBFbg3XfeA/DAy/MDL48LORVrjB6iP82l7PE4dOf+nFy/d94+8dlnn2OGBOXC9pm1lAPP+4TuePX+pZC/Ps/jD6QUe/Os87Zmt0OHmth2kqHnEKCiXw3UOM/7Nh6tIxWW1suoii66zs2ZM5h0fQB2BJv7hJFKR3tS571OGfCRkj+tE9x9Hl/LIMe89wvO821kbrn3yE9/eE7mlUcAyk9qC1Faixqu8xbgAiI25F0BPRT96qRCGRNrq9jRCjgm7JJntNJq1CBEkp1oGrICgUY1y2gDKNI2kVgZbphEjU+3geOSq9OpugOFkA1GWpgYaXE3rvpcvP4O7zkUpiMTYT6lLTYjLznnKUc+CxVxOAvR1wccYq6ITaIhNNclrPiJcBKV3vv5j5/N6bRVRFYtBLMRC8VEndNCQi8Ma9Hu4OuMSCTwox/5jFtofmgbX8XZKBdJS0pXwAofTRpS5haimtb2GBhxUhSHKLmvz2dB7jpSgGvXsrFoLIN5FH24MtGyzbOiB76mzAoCq3rEpjMvpyHkfFChuYlwK5u28DJ0VKBZYyyQt6rJclZTp5orX5sKNjf7iboBs489PIRKGk9qP0QcOPd+FGcxTuQWwmhB5yYWJOTnSuIacl+KGtTnyzcm4WMuZCQ5BbPMWljT16TeAAAgAElEQVSC2WljIXrhmFUnsrXPLlECEiHYRBsNUXc6SoJE+X89GbpHWNC9gNB8rGUuoy7jDTe8MtpLkDNBMLltQleAbkrJXuo9RpRYEMy5YIKMSeQW2FWb2RCWwn0h9ti4hOI93yUkfJhdc7UD1/WCqvQ93Ycz7Y8jRy+m9PtU0rVZVvNSzBZMsGN1Nsl4G4fgOOcpbkbrNrt6zC10dKtViahQqxTPRED17527635wvwcR4IgYGe7D418HUlGhgWyFjPpVIZBxbSINVEY0o4tAN53CdLVQijzRXbYsn4pStOGgguR5Kby2x5GIMOLSnPUzZjAilwOZ7EZ8ALBxHuvMyKeGYuVrTcjD2o5MD6w24N1vZ86DDvslKhgEHo+TqyYmT8h89GG8qYeIXO13mkBbrZ3pg6OtDfkMI4JXkEsWwVl0tTHLqjvqkqAPW/fkAtO3GyhD2rlHlpeUkqHfARZmLFpd8UKdNt2hY861FEYLiwT/1TOlsl/J6awOa4bWopRCK0POE6/TyCLhhB2SfrEOHNkZoGTme/MIUoPt8jplvxWtoXpqLEIkLQ91L/MHPIzH9QiOQJTidzu/TRKuUQIjD7i5zK6UHixJVU+Oe0ebfSJSrqk2cx+UxGvfonokKHt9pIvo6nF8Wu+e42D0rRATnzXWE3ysQOhvdXMHXd3T92h5gVa1/k8XNpGDs+DYHOad+4AJYVNJxeI+nq0pVi5DtjZUMdrdp9Oy72czlIYnhKMxn4CyNOWIdQOY9QIkpkxeoRaBA6GNJtSX0PKP8yVo3et3LsRINJHfmzpk2dfpz69jHIbUCThxgL08IvxctffX+HsqCkeKbsU/MLzl9TgnJkP53PVn1jLMuZux/wEBPVdUoGshnt50yjGt9wifjWu9/63/dGzoHArZ5CgWOZiuPenxvvPzvzzW2JbahHMrqEnK6d/cY7735HkU9Yr5HfJVobn3bCy4H+yUkxiywE23boZRPTyW+0VQWd3lxoVYvI/HwnW/q3l/nmjHSJBut1CDyE+MOWIjKf5+2WjoWgPpDr6D62pClTVCRPhhI3KTLeqGGvkJehyZSDwqiUeWabD6mBatJ7stUJ0RWrBx4bTAwTFbh5XyNqiIyZy7wCxzK3GlhOQqDmJv98mgpLEohtYuAoyIiFzqe/EQ4bBJrPeymv9Wt+sX2OcN3ycrWuP0XiuxvV/u2ryfMY4nKdTkZsAIscWBiNS8qtEx52ed2B2K5fWJIMqCQG4WLUUm8NbP/Tq+8Cu/ipdPv4f11nv40f/zv+BHf/JRW+keI49IPD/E21/9Wfzw99hLlG5l4u2vfR2f/8m/w75e8DN/9b/Dd//nv4N8+gKe3t74/JPvAfEW3v3FP4sf/tv/U+td4bbDMsNr9g/D9CVzJid10FPaje1J4I7TvEX3H81x3Zr2CstbyO8OYslCKTKlNev9kIFEkAR2AVq5f9lTdyn7Vgde8d5KDjT3VJ/p8OS2Oz4b5nBOJoGqeRLySL1XbksvV4eGK3n6UkCg9unYv1TW4fvuvO9tFoFK0eZGdui0f0hqUbu3dh4TJogsWF0TcXQXp309mgSiEFSocGFGFaKyI4FhjTsddS0trfpQILAjm7Sp7xAGF9HW6chpS0aflddW/4l0BmLtcwtthbhwU/o8KAgYnEePrbwmjmMJojLcuYmQtt0kXoGhumzUItjoW6iQjwcOba2J5448z0o3QanrH/jib/xlfPwP/y6u66H7n+98iHz8GPloEvO9D3F99inOL/0C9vf+CE/vfhk4Ey/f+xhxvI23fu5X8MHXv4L948/w+MGn+N4/+/uIpy/gw1/7LeR3fhv7OZFvfRX7+x/1ugNPH34F2M+4PvuBrNsihwK6Jq4I5jMd642UINDFWU2whvgLb39yOkayXCK6CpBycX1GSOZe65AAayIAhrPFKcy1zwA2XQmMzzEC1C6SqrRbPmOQ6kKr5ZoLcbR1n4dCobmgiV48ZrsTESd2FLm5Y6BXukNSSPsmR0DKlZQARmLF020eAysX89/lW3P6Y+ant6ASdo//qImjHzZ6AQS6CHFaecRYzHk+CGeA1BSX5zUsmu7RXO0JRalIGMalBvAEsscCP0OI6gkeTzg2Zgsvn0t+7Nbz14hsrbSBAZD7uIWheU9MF+sn53d1cxbA/SDRFnIqDkHOOODW83WvD3/zr+Pp7dqUcb6PL//l30LEwpuvfR3rvZ/Hh9/+S3j/1/4avvTt38R6ehvv/4W/hHz+HG8+/CLOD38BX/gLv4H19gd47+u/BDx9gPOdd/HW1/4cnv/4/0OsJ3zxP/tv8P4v/Sq++F/8Tbz9s1/yc3M95fbBgq91vno+G4vclDY070K2kpdomeFc+Su2ivlKnrfWRuOC6440Z1EbcsoCN65kRp+blKqJeMq298cIG3cfzVn0KJnr/1a8uj9lSpwSZf+nyAI/L01wj9TMPRrtknm9vF97j8SawlsXWEPo5lK7CQhgcnDG/rmhXgu8ClrmA8hdSKGF+XNPXDJJytfuWZa4CdpMx70dGiPiMrvHwoSw7R+r/T4XkP+eSTRWPFJ4eBWau0364FH0fr76/E8RePnHTuslqC+dR1JWs6/PfPLP/yd8+bf+W7z/Z7+ptT3efRvXjyqz8/jCz+H67h8iEHjnz3wT+9M/wCf//B/hu//kH+Dp578FPP8A+7NP8Olv/zP86A9+H09f+UW8fPT7uL737/HyyR/hB7/7L/Dy3Y/x1he/gM+/+zHe/Y9+C9cf/K/43v/xj/H5n37UJ933+JFawxV+4qncSGCjERuJZr8Wng9dF3p258AElKg17yH317kySLuD4mGGW1PJgbPGZV7H/El9xTlJXMeZa8HPhQyVnzloYQein/IjRaKCymGIKSu4535oL0tR3D/PPcizXXS0h5QTxutl7c8ib143AmEYqPy7WMet7HfFwh5WM0WsTP3X8IswXz4TBMO0mLp3fUpuRkTrrI55Y0v7zYOMRTRiJDlFasqQectfCAAH8xsigGGl0RYoAZ1tWhWrR8ejQ0x3oGpM0Ez9fSkwjhsoQWQItuZhS0jqM/X0io6IM+k1wLShoedYcSjqEC1QmRvXx/8G3/mH/w7v/eZ/hS99+EV877f/bxx4rjwVAG/9/Dfx/Mf/GwDg6e3ER7/zfyHiCet4C7iegQTOt59w/bg4nrd+5sv47F9+jHjrq4jnP9Vznm+f2C/A+9/8Nq7vvI83X/9P8PjT/xef/cl3tanrWeq+zrSFeBgZDwRi9EGh4eLz0iD4J26K1MVRC4CNyRrordZxhM47TO37eB/QemdJe2/WlJthziV0/7rnNIyUlWWZo8FZADD6b9akDAVT19m4oIxUcoxEtHHP8iWCQsumEtuSCucVAhUiciJlm3hEZEVx+vWTGnL3wFLWd8bQCe2ZnfgCkAgh895dqJTOnNChryn/Ej1RDhU5y2++P8jQW2cr1D3XK8VGTd4pyD6RqywZ/WNocw4tnM5FEDxsP3Ge1J4gfB2WQveFjxsgWgI3fH/yxlLjdo2ZSWeUVn7+itNWTMJLGEuENCMEPa79QMaFT//FP8JX/9rfwPrDH+Px8b/W/d/7xW/i49/9H4HjA+DxiaqD3/zCr+D5j34PWO8h8od9KPDC+c4bPD77MZ6+8Rfx+b//VzXm40Pg+j4yA/nZH+Hjf/z3xEmIfxhepJPP7F/olK+WIwsC16KbIXFuWqky6qQir16f5BxlhehJBBPPCHHe2uBzfOlxaK75Jl2GgSpI8iObWqh6oySKuhkkI/hSMJ1B/GozO39izNn4fZZdgDIpDqjzdIiebtGPBPOjgo2tct7Dsr/z0TxYWjcgseQqjP9oEXx2Buv7B4mX7q1oH8vNViKi+ynQOvbrWZSOD/ulHhjcR426XkvACU2pTadzJdJwXt7d4Bb0Pi1v8tqc7hifg08vS3g8ukd4vANy3j43EoT4XHy9Z0jvTbcNHJcg8z0lOMZ3Fub47K7w+d/62W9grQNrvcEHv/5X8PxvfwfHO+8CfZTkB3/xr+PNWxf284Wnr/4Snt5/H8fTifODn8OHv/xN/OB3fwfx9s8gXn7Q/RreQeAFgYWnD76C/NEPcawD51d/CddHv4/AhcR7ePtLX8KKA+cHX8QML/rvEeKkZbz5zz3PXAe+nhRkSGb4AteqJ9CNo2/3npZ0w70qxtryfuKg6jper7iNx/OfN5kqJNOIW6d/MTzKsGiN1YAf2kdLiYI2ZjxNjnOkMYRdi2oMXM9glNn7tPfuAlEFhEDmH4/d+5+6ISJwfPUr3/pbkU9d8y1V0wbSDzkt5eQX9ABivDlIwuscTTjGPcYEaTLBzQpd06gzZP1vvisAVciiPl/t28YCDgEgalnrBM+AwCCkAkxuMQylssm8tJhTqc0cjNV9H2YkQPkVgsrRoGSST2g/lpu/UNySgobGd4/xHx5jv/fma9/CB7/2n+Pdb3wLjz/+bfzw934X16cf4c3X/2O8+40/j8//zf+O5+98jMd3P8LTB1/GZ7/3L/HBb/wVvPnSh/jkn/4PyJcNvHyK42u/inf/zFfx+Xc+QTw+wfMnH+P69Dt479v/JdbxgnwsPD76V9gvGz/+w3+N93/jr+Ldb/wy8KNP8Pj0+0JMM1+B8gDK04TvfK5EhSk5b6+UInKmJIfWk2vhPJHoo/5GYSEW0Ghpd8EZolH1QMraqL3poxdoVskmHBUxV7a9ZszNyMo50r6Z98CUgXvIl+41uKfCijPm/wfhy0xju2v3PRz6mmWaW5I8EbIU6ix5AJ5f4te//V9/P/fbH6i5SU9a+eCrQ0Do3AKnUHMy6gDgrc+yYxChH2EsYRGhDXtj8vfNvIQ5IYoVu7aCfMrrwqna4DMUW7CcPER2rQrdpJnUJVDcfu2+ngGSP4AERPkD040aioM5A0iATW3WrWBpvXqW7Bz9tDCqKVArH/ZDGJEXaY72dW/E1pi/Ob9KYpKQWWnXpSofhi6mnon3FdxuKK2qYYaOQ+OE7tT3VEZutDzURr86T2CS2XNYLLgqlzLvY5oVy5gZi3XfPTYd56KU0AGe8zFzWo51an2ci1BzyULCqsh8uOdlK/0593Xtcygojpk5QKMQLE7Mg6oos/4dmvPJ0WkfUJFwvmbBYzir1U15oHvdCxindCR2XjjWGwCJ63pujub7PzgrZfYNoHzwS8JAv64U/IWk5iMJtQEnJrV2rWFDhn2gFAuRhZ2bIcBCGhagbVmhBLrsGqC1JbGUaFKQkxLchKPcPjpXQ2nYzWXIcvG6R++/12GnUhyld6q/x82ih6tLGXqtz3QKfQyLJ3/ex+VZgS7sMJPPPV/KJHHb4jcLQ+LQQsHeHMBuRVO/zyY9Us69ATNDAofwZidBee91sFW0VfuQDVtm0Rx5HUaiiJLmGnj+nTtR31u3M1tcXkBlz9yT6eKQK1ncvP2sVY3pOV5xFPel9TPRLmTTE6yIX8syj4WwIphIfElmRe7GwnVdOJorcHJdu0hai5GkHrUnqChyrLWicRhJkjfp6DlNJytWtXZXp4J83zXG3+Ruv7/3C8RnVnlDnAXHQ/CZgkNorf4F0j2DE4hiTN2jYam+pDZfIHHYYulxbYkoJK50pZUhGjEZVl9x+JTfd+EZbu9xEaUzB+Goe2uTO+PNEH/1Qr/OGPVCineYKGPyNkFmPnQ/jsmp7FPYZ7evul+x2qk5JsKDMKXzRRjZOY4DJJdv7PqwhlVBjEZAFbmhBSu097h/nsIc0cVFdg+yx8k2frM7GT8ZcWB13UFlnbLSGf/BH7uDoyPYWB+Pi/N+V6K0qpPEq3ndA3T097JUlF1fhsnrmY914rqmvNHdkUTc1r7mcc79QuLS58e37mOQMVza8PP5ZCwRt+5wctvT+UWsGN39bEQ3NHL3A7xD36Fbd+3n7s4fOE2kzPizpqona2tj1Dx3/wQSNihXIffGhrtPZQ9mX88DNjUkk69HBhitBTfIeBM6Mmy2xXxPSBzw2RZ9a90rwYY0pdH70ejT9u/RY+KCJDfmIKR4slP2NXNdnp/LkC6xtWGIzqrnYrZxup+JMuwFcjRkYUo5VjcDImTeDzD9eW+2NXTH9KkNb1EfKkxZQxqEQhwFnwsFlJVhirrXfW4eH6XQe5jQuVGQ2ry11St5qfqGHSMSNfqixDBKSmtO+HduuKzFq8Y+zBge52oojduhSikNko6NYGxE1qtnjDFGDFkHyDnMaCHnu9LAa97WQD913U5Rp7sBRuqGK9IyhCa5jQSsEJXGEF4HtdqDUV+04daTSea8T+Z+IWK79kPjLLhRc3iW/3i+0i7uOpW9FGtmhktCWqvryDfzGUko392mCuK0NkyjE/IKnMByAwhfqcVTJNPe1yiMitLUOJE7C8L3eOdhQnPDb7lZ1w3NJBpB9YblOAIFzY/u3ShFtcdEj0ItpOPVaKQyPx/aCCY6TXhNV63EBl0BKQZ8Wur+T67cIAuhT/X60AoPX39+Cp3w01ChPxtaB72GKnuuQrvoJd6KhjJpiDDcsHqGR+FxDrdvQvHsY/zot3MtnZJNzc+WCrWJjuVr3e4zolQVYpzGMJDRcqEuXtMtSTCAuF+565PH2+zw1vIwz86pywyDkdlFzVZKoCvT+8KRnG3xoLKW2r+jxkpoI081unS3e1xGMnoNWfE80WaNSHzKIupZeZamvdS9uZ8G7uHXkHRkQhbZY59to5KCnP3YzzYUytLTQgKoME4LUwCqG6mniH4++8HCI+I66udYZyseWzJl1pKbiMAxeAlaE5KwIurIWvcmZSIVN8jeaLa+z7KEYR/nK3uBy4c9cedtuhUh5ynGgpL3kLXtJxwNhr0OSwIE6Ct+XgoR5xZQXH8TQbQyKgVZvT/IFcBXvRkH5eCA5CJdQ+DaDwR7RST7KRx6rrK4Z2O0qSSp9NrdvdUDhRRw2aJuo9BFj8qEbBmupMG68hJMJ5Fst6LOCA1dT4VXfE6Nbo9N1MSh1qgAOuUr20IfPBe1rTUWyfZE7lEpG+gTw7jZLft89llFC6mA3ps6xCiECPjjHdeu/iDHh0RAyhhVg2RUk9BpdNg4E30oQ7KxqCE8uOCCi7RchHYOI2byYUfF5CDPAmFGn/NB7T8fbzxsvTeVl1/lDzMCfRzbcFHSm43KjZl3r+46BOrSSdi3DNQ+ICmJQuTzep5qTu5ZenMz1OcSswqQC1cwGv4MyFH09wd0Th3C6ycgQTo3BufhdbSAB+zsbYWN6XKpaZBD4RwXmw3PBCNo3fmofuYZ1uNc64OcH6IOwXl+kugAQCMaHra9u7R/ab0H+Yqy3uShdl59li8aMZTi3/lS/FqOhi89rol2HP2C5rA21igWGwq45PIaKQbZyYQz7G7DKcMCGrJWqm30ciB9/ljB0fUg6Y4hK5BMcqxlHEYiGd2asEQR4StJLQp3nwuRKgEGi1GmS8LNzgnckgUbMcJHQ2X7q653I2zmgES0wKFZZMpqM1xZizsgr1h0enIpoZ7hVMEzbSLgiBMJ+vrc6JUpWVq6tD8QDrMRdWCEIXvjznvcBEAW14sr1iABkrox3wu+noKsXIpSco3EFlDdye2zTySB6bvCdmgqauDQc1KpTbKW6zifoXS580cACth0oRLMY/CYauO75J8QmuPty0+5opUPIi6SyLWOa6Tua3BCaD5kp945dANKC7jZmgtS/89GpHrucA9WPi+raHnIEHq8R39nDSKaz8pco3rcWl8fe7goJD1Ph3iG1Ui2Nv3dMNWccH6YwsAyjbo3Sf5oIxUan3+q3KM/D2DlkBd1Bk+cNAS1IXJYinrt6jMxd15j8wfYgYk5BAUDVzP3zGWgwDIph9LQvYKICHoyHXo69HosJ98wKct5A4Zm02feOqbNIUpbP5NrttwWuAhbFbLbZPonI1/McmrMMweCAsmaDZ8kX5C8WslfMNQkRPYG02f6/eICqlyem8aKInR/N2913ch8PoBNXV14VbJTG2Y/XqpDeUT54HB4uxT5TEvndz23SVmQ4qagtzK9zbkhv1Ape4YKXRAFVHuDFU9CAZZ53qsU7t7OcaALc6ynkb7PqFTg4tGMGvfdUHJ8c56nEZzXMrVD14hyTzcCQxaaX+j3zYG4R+ncE3NcDhd7LYo75F4q0toFeeQy0NwLwBygkjfen9Euj0nEJxZOZLsha3QT7s1WBSyoTbC3ejZKs/WgN8nD/ShYKHge/fuMWkDfZUWfNjO12zhV3S7NyInfW9dUCKkXlwkvdR83LWFSFq1uoRbWsbSFUs9JyUkLRP8ve2PvC7d29pEAe4IWPKjXE4L2ZcwIu0f+vuBfAmOz8X6as6x1qOZEJNRYV9CRgHXgerzclWBuAKNZcADX9SKlRwWSmX2maqOH6GzFjMEj0ZjU0QnH8dTPtKFmIP39/tQNzWjuormo4Q5mu3oY36OsMIKRmdX4KFPPXJtqRCr05G1t20qWfFauAzJbnlty5P4xo5fym2Mc3pyRnr4A9I8Ak/+g6NLY4jeSe++HUNN9H6Tknihu3uMWVgfD991wqiN/XJu9y806upG15Hg5D8P1MHxmyP0kZ1GaaeNcayX21D4tqNHAuzftWnZJ3H7d5FHEUYNCuQw8N4Hx+BLIkDYjUQp2iSb0HoJlGEy/uTdQrGaMIWuuJRnWTAJ642EMz6miwO7G+trQFqg8CfvEhzbAFFB32/bXvVFoNWcWXTesgcelNu5UgiTHWnBXnMiuwHWv1OECxInjcASJ95m9SgAiji2kw6ZE1XCGMzMjHqXopzU9uumurSerRxsdjlO5JNRxDOQ2nw+wYqFrd4fKdFmtYJmzsIzmWvg9fx1lS47L88r58CblWjO7uHXSRFEDqVjuHcaOMDpxJXcj1IH+EkSYU5EaYfJ5jQC9btUlzjkUvS37noe+x7GFnq8VTwTucnnfcwxxE1GI10LgzCzNfRz39FcyvnQj1OVqJzJ4WA55Btb9V2UqTyPbY1IpWLNLdOIq7bkgBSVYhRBkKiBSNo3p39J+yqNgVuKY2LbWaHcpjidw42lTtoVKlrQXxJDApjqD90BghYlGDkU4Drh/s6BtJWYei67F0G+Nf3c3bs4pAOx8UWZmZdVdLJh2angrMrZ1U4s6knft304CtBSgbLA4kdsZtFyWOe5pCYeikuVri5r7kgvE8ed+1BjpWpJM7fnIsTEk0Fw/uY/2rWtsKZlibsoe62TU5rnd+1FuCbKnr8fQmn7ni46RuJP4bG/I13yPJX6t3iFpyamZ9RqMNES4PZ/C7eBwSx68DlvHTzLvCcG/y+XWc+XWOvI1nulzU3Qy4kbJHIDyffaF4+BxHLvbyJPd7hx27Zt+z2E9P9MtCiEmvSE3CEuzb375z37ouoyspAa4e8Euf2ZozxIFk0JrucDGvuBwlXpRhZhgwgk9VnMpA21oLNB1SqAfY77md2hBcHtdFlTX7E02YGxFX6D3s59RBCg2dj4krHxNnZbgZ9U6SnC3noXNgW8FQuP7WoP0RqAS10OmobGT6TwXCCrQS88+n4f3YM/Iij41csMcy4YOvqab1b9zPYOf6zVcw6ILmwyox3/X2lNJ9fpTxijcQYLXSk0yQIPDJCu9N67FuWhCVnuJCqgJ3LmHqPi4ZnYVtvYB51bzNtZdSv8mC6m1mL/fvp/7Nj5/1smSAeBcayGyj5tfDpdRITOuzNOefOpYXfyIo3r/RTXEYU7+Ro66iIa3A7YKOo4Fo6WvIoy2Dkg9SGDhCPetpI2hgqhFYYJV6D5u1oPuz0kUIZum56wXin8g455BAN5cB7NFI1wSzQOh4esztEdREjvfadEE3DOywGvP8QUC0QV6zJkot4bQcev6icTBkK/W47htCCQAnQRXU51x1Nwuw+sQkchwZCqpa6cTsGakACKoO+rDjdH1JhFwEtsk7jIxjwxYsXCFLSCfc/G0L82b+Sr+zHNSyg5b0hYCm1B8uL2sFFUjoZvrxsrpaKmo55SsUTfQDZGcY1hwaN2u/YAb8qBl5JLbsBBde+I1JBrTgUNj/0ge2hW5rksyhXZDlnV58zYO965G3DkUGKOGe1EHnF2503PGY/vqJhTZqOSXhAiaCelAv05ucoAHyoBTxDDYWFimRO9xHYiH4PWINrqoSKSWJyEzPb70A88/jOFPocrmVOo+TT71dcimO3t069oMMzovoNnpPtX79jq3PUk2WXP/LTj/U+cRHgfnL2W+xxzlWBvfm/fXova16b5VlqR92JkOPPmYHN/jPfVGJnLnaIQ8ZGM8q7gErctPXs+cVbm7kxS0hS1p8OdzXHt7PpIycc/bqfW8ND71VRlrubPnZve8UkY433tLJny/Hhfd7W0i9rYeSZ09ZJ4yNaI4uVPPmlrX8XmtM6e55ajHe+P/2Kmf19sMNIT/vT0HNbZtOUPtiTP3DrLGHJUsLyYz6nMr5eerliEbJtN/by5gm8coFTiEGlXjH1oAdkRy0ojgbnfH4uDZafwn8hQSIqB6ZjTBAYIVhs4AHUYsUhRSQvV5IiBI42a/XmW7s0DJGaF26erGPtsyPceDZBXcH88yk6mKc1FyTFmi18pY14GsHZ9HEZ62Sps+L+iHc919jR4YxF8p6Q19P/I6TSIGBbUEMUd0hG5hDXmD+QEqZw+2GOjuUagwntbxplTbldkU6IXbEw/Oi5uSbg83EfmSaBlCrynn6bj1a6FRIrdQ63gr5kLJ0LUvWB6JFBNgeveeFd0jL6a1BpPI6KIFDs1BoWXmfphrE5KlgppcD4zgbiR/X6+WesyvECRT1bnXa5xnxIpiVUmy9CYVBPYiVQ5DZwqqL2ad41gpvCHY5aSSU5PN3AROUJFCM9qSEtz5QwbXTDG1JGhwcSt4uikNAJGK6kx4miBSGGobdIdScLk2LXBtJ4TtSQRyI3KcIqBqIyw47GshsTuB3A0vmX9Sm5CCWrT+/jYAACAASURBVBdaPiphKq4IKVjm88eYv90KNUbiTa1Dn/I1NlTNm2H/ZppzhAS3ttelk+PaNoEVxmTfg5sp2oFrBDP4f8iVQ6gPCgAsnEAAFzeXxgnJ5k3B6ylmxIluHsnIOve1lCU3B0AXNPs+pVToHpVqZvsDkuugLIa/c0uRT8q+o1WVafxUr69Kix8S3rIQFHi7QuloH2W6omFQVJK1XHsRrV1dPRxgvRZdxt0ENJsH7XShZaISy67N4yNaJmOV1Bgkc0yGrXJEYmbs1QQdcWhTSqDCrd08WU0ULcf6AR56O6CS7sX6jFZYwzL5+6HrssRWGpaTTgsyFIChIEkqHzPHsBtgLUtBJWwuvxZWDPA9RISlTxHTqOSCMYuPhJJRgYR6CMZ9bnsucrYzLH/W2YGvFd9Q/olxn3p5gS5IcwCj6fB0Yjg/HI86TLdin+s0E+DmE9PnZzKQ1lhCyTH7/vTr76nOIwoR8zXLhDGF5UqfyTvqoDyTxF8Y0Su5ET2mMIYp/gtee8mjCe2KaLzc1pfy5Uxpr5HmU/fj2o991p9z1zg0j+fnXeP+3gM/Ra5jRMiA2++3+/X/zxWRXNLsGyUFtB/fmrst3Cj4AboXgnLkeRIzU18Pbfb6fmAunolKWuHW9gCKAGvr1l2vK19oaXxHnI10SDzFbYJI7u1e4aDFhiG0n2v1BG6pmNXEES9JbWvizq4Cld2MLhRqApgAE+vUdeZiJS2+xD+xd/elQDRBe3S3LmZr9jmxYEEbUYh00E/mqfRzZfB+vQJhkprjmOulfA8pbnRn81bOHNNtLg6NgcV6DDnz+rcjIAwf+K6tv1KzbVCMOGioLJOpsVtBirjF1nWodFgsScs90SerpEveDujEuLAxrUkvV4URDuYe1fx0XlEm1nL1queZBYjOUvb8t9sZxJ7QWiacI2SFwb23wGpZZmHaHYFylRSt66uIAFgLy8FInNd+xEEfkX5sbyzGiw2HVvMHVZdwBDPHrvZxKjYcYDIXy4ZPLUqVhtt67s4SrMne/h6yewhcdawgJygT2Nft+sExwFV49vVcBbrzpe6BrepF50FkR2zcL4DPlLq1F2hJsO3/TWSAbJ985UisSeTlgrWIhR3T1elo03K6eZ1q3p/vfhO5H3XPdhvILaBfw1AUF3Mvhs9K/zYxcz9Gp/Agn0HX5FUrQZbnq0w/tYG1CcZGJDHI7kuKJOTGRS6gN74IbzVVQstmn/OSqPFp3oi6dkUZlO5OH9w5OLtT5GsM5mhKsWwpvFIQS5mrez9wRPMPSMspjIfY+xI4NI/ReRCq2jYx1vLKMfTLKzVne28lZa1V7h3yqq3fipI1Kow4TlIyeUTmvrqyFmD4HC2rW4iNqQoYyIPnoTb3gY3ziKPK1tcBVmwGXOteg2vL3ZltxzqxNq1oVigGgYhTAnn0QNbRmWqdKLT3vZ9lZXkuTU6wt2HrN4Ws+BBtZZgHX2/ZYtUp5f2w4eu4p+hGdOEYU5RpWaWhZeDrmYSCVMjjxrylrBaOY7Zor3GVpVvVE0AMPjNgR8u40Rq/6jI6o1XH0C1k+tBeKhLiPv5wfdQvNbc4I/Ig1CRWdvAzdQ0GUAV3V9dj0OdlSTnvo5J+QGOpczXcJ4FWN2NsGqLOgXh0hAAM46smyfUuXGvD6TUQQmKt1JiSiA/R1hqabxuJ1Nxrzge8UQ7Eemo5JaqqFPO52BELPAHulr3aYziPewSn6qg6A5rh4HBx3zp6XMwjihaqVnjqZZpEjmEjnMyeZmsAc0kLoftynLq3VtIVsxeVFg6sWVY7/VMnd8CWl5GP/cC1HyBDXrkX9SCMJNDfY0LJli9v/7B+OiGl4e3e0+en5mdatKEWH8sJTznu7e/7OvbR6KZwQlY3ftG1kxvq3rzlfk/oeYhwMLcumVeShPUi7n5qEYbkOvR9RkfIgezrdj4Ix7iVnPPQPZVIAypCsuZWFFOpTZfNYyLyg9ZdBC0RzN56fe+H5GWy9DGuH5h1Oxdmoljdq9dQY4dlJq2kJx9Uf5dFDUL3IQ/1/p0Hqfsz4cq5NWqBjzKcUhSaC193chQaOxxexxizxiCupI0X3VrEeCbyY4yG9If03LU/vJcoD43A90PzvyLgA5rv82dQnGNdB5czI3NDN5wromPN4+Fi2XUArd/RvmfDnz7JqbR9i0UclfTCzbjoB2Js0pCvx89Guzcks5zQwk9xckPFbAsmiPg92edgjoQ3twSRpBkITzlv25xF11ysWLiQgxzs74+oDIV1dquq5amNWhb6RWOQgI9TrMcT1dzRFwY5naXy570fWMcTgvUdEmfY9yY5F9xIFkhdm9xDz+sEGlJsN6XqkHrJg8UwyPeAJOnw4+GNvdbq5jhck+Gz377j+7CmA+SLhCzoNo8q5F7jSqJ7FX6f8xzks1gIGVAWastCQLEpINgrxMlW89n66RBdYUa38daiAO4qn5ns24NMV1xjjFRGicQx7xKOTtAti85aJZ3BWg7uR++fkl+R9uMAZfV05TMOPggd+TkpBMzookDPAhamhZIA4galADKrc7cvyO9gpyc4AfrIijx0tSC15cI4XbsFiL7y3o6D7xh+ZYeJDG/Ln6Q/WHPIgiJbwwzH8bMLxbDob5KBhHzLhd6c9AuVlj44CJSkitnIjS23gFp9gYVpW0ijhINpz1QShNssz0a/zh4fhLBagwU9kxqzZN7ITKQ3XAkCRdTWz2FeaPNM1DQJWSPEsk6ShZ1d8Xi6uQotbiMWbrprv0wVAboJtZE3riHA9MVZUbmQeKjV3b4pkehcjc26IbT3nVdxEM39cL71rInKVO012LmB5k+qk9h0M4oPWJxrGPHlnnNY3ILmKa/hFY5cEE9myU+yCU5zGXkBWz5Aj60N5HaGK/dQ7aufliIw1mDIgmVbd6DOxbkzcWS20PGCtNhL1aOs8AsKHHVdLJzHU6ERhM6BXDhGh2eik5FvAT58h3oG4xwg001YRE6l/mNCTPnAPRblEVgTU7lQiXAzUBEsGCHRpWI/DNm74CTum6XQGEArQAp2aGSU0MXFQ1v6/eiYf5p85caJcBEcE5VmToVOhgOw1pM2ELkFjsHhRqd+O509xz1b0EA4O0LRKn4jkppVnI5IKZcjAsdyNeVJN2/Z3bu6IDEQ+v1QJ6fQfYQgwN8JidunXyfQZ8XUnK1CCL2yTlgCGFXpGR6Eqh1VpZPHvN+SK3YPJdqNIafCmajGNavyZthXAoFLHMEl2StZ1CoMhAG2Ohkh1rj/u5Hj6tcQgWNZqTji0QiteQkTmY4oUSl677QUNQIhF3MiM25asDU/qCnzKgSwr2oUgi6lJmzPjcf13CXL0CRnW2iGD93oNBHdkyD3rojH9r+LjbbroEVvBAIAuepBkguJ7F4UKOgN11gkEvsy2RTRlXQrOrt7I9rfXH0c2hQ0+uZYRF29mIst+ojurBSnH7jx0Dxmi646TKORiwi7yn6kBYq+v6BjWJUjgQvV/s8FTfbJy5KOLL9Alzej18lCsxONQHodMrEDsPWkEnKWrVvu9fm3naR3Xc9ScO5s3dda9Mcpa0QwvdbwWlflKn3uVl7bjXHyYuSm3t+DJFbGZGOJGi/vVDK11sEJru9ftLYmYLUXshK1iPxYPJb9+dy16Xluyu7Dt4Id3ftZ99XHYZDXWV7XXnjfPxMZ10DgeVNcs2Ncdr+KzYOcLp6ch66uJmJqORRhwsjR1j5FdqtKAtGsVPAdj9II5CXqb5XK9J/20Zs0ifZ5QaKEkC/tnkDC35MpwmdYrwFrA36P6Iabi2PL3G21emJFum1tCtCq56VkoAGSe7JnTYuPD5hjmG3fy0+mRRnZgbmVlMPnC7y+pv9gPJv/eMwCljdfN7libRkpaH4dnbEpRCOkWYq3wXw9R8slfX9aUaoCEXfhpJ/ykb3uikJRNsazSrnIbUkZFP6tZCcONDkPwC3AIIWdyD6FnmO09STy5EbYmh+7OSRb3a9T99VnpvxhvMZp3lqX6DHweXl//n6Tda7PQDVcRskQ5RlUlv1ZcVw2JJLZqOep1fIzx5AJ3iZuz+q/Kc8z8Y2ohfuec7CiNMK54sARb5TYhH5gHTrUbf7rS91ePBawnvSdA1mQGITxD2S7Dtj12iNct+9FGXBJaAJgD0P57cifiJ8r03P0IQxNjwUq+9r0yQsKP4NJWNLc+tyUl5Sw1FWdThxAQcWdEtzUIrTnl1uQlL0M7dZMGGyLcSxXcAbnSxD5aBTjlOyCuA8cUQ2IYvjFtBgLpyIFLYniPZgTEX39ikY2RF5PEtyFUCi3Tq+r+QCNQ4fpWAawRm4NQ3+zt2TdWzgJIGGObDfxDvcpCxnTEG0w6Y4EOGX8oOuG4nzA9RHX1u5go0NvaED8Xb8x7weMmhb+vxUpOSivKg1r6vsVzqRSphqbZLc/H2upARnDwJVWTvkv51bNenYAEVh5qL4lV1eZdhu0Y519wlkrzwhAxym2vDF839dir9E+DGQLChre7PGgJAV5khSPQeOzOQS2geYStsjCCS/vm8N/A/aR9gyVShBsWQT1h//sH7P+9rfpK3jBGS/newVplza0Q1PtK0eIQ7DvynV3ohHHrLGjiCdHEOhitIIZgsp5mQRTWXPASTf9OSIahObx9XF0DvHWNyzkNgoxrkWGPUo6FaECOsciqfOYqMM+oonFDYAuPtzOzi0F/fIaOgwF2BZvHD7kg4UGUR3Gi+IzqOD5PzX2bYIzqTKCt52TPTZy75t05KPvBEhWaw4qqvNSdxAiD3dvu60eetMl6OJOvkT7DDRG41BjyfdYM1iqeYfs4rxJUrMTWiH7up46bxHJxFaCFtffMkgOyXJxZu6YLCwfxt2va9qZaRl6iEs+z2tYSXa7CBwzxIfcCSf/FJw6cOUzDhGPZKcJ7Ut45J+DRWnW3BNd2KcD2CFqK5+jk8VIvqYX9S6IHYYEIBjdlh2y9o+2uCFhNgFIpcZmv6GNJeQDH/fIkKesD4DragvOrEOQIAZIPgPkJoxaePaHkEVHJyRc+Wg+AV1MVuPnkYI7L6wiMipZbiIAtAC2AeAZolMJMxRXSMBKZyomA11GI8ZOuG3QdkM7ojKtMpW/CL0B5ycK3pSl4NkzJoLRc8m5WVRYuHdnDyzEMgfgA3pmqj1J+bbw0WnuvTUmkgWsXDh3suyd1s85WnHeCs+854o7OnD2Wna7/2RGdnQ0r167rs5ziTJgaLlk5zOm+lMxUtZrAuoqtfH6GeznTDSQ3aSUmquv0TCbk4ltlnwik5ANoLAaRTDN94jDk560qLbhVFI81AeZUl4az6a18b9lPZL59v2MCfVgUH7HzeIGV/L2N9v4oze7hHTyHOh774HOmuOomNHd0k1BWz2PNd4OOXefg8g5f1vXsRJvoeT8cL73vv2btreqgkzmzbm/RwumkEp2NH5QXrhuWGDFkXJU6Ibx9DqORohgJnOxhoOM/n1sNCJGXB6/nk7jgb6rfhF9n0Py1g1mxjWYY+F5SD1Dai7RiAqSL8tbj6nHMHktqFdF3WeNcdzl/o4+FlppYri76XXxfoghq15D6eFthEk3R/N+k/sc/wZWWaOG9Lwg5mD9OzdqwtrYyqZgFgdkrczFG3B/Crrem+E8hzhVDzDw3cQBt00qmEeW/aYbRxakxF+Kq6IejlJogRFj4jjb/N5Wo5y5yEi7IlIy/TyKImgRU/OvZw8vGJGS0oTR5caicNHW2olvqkjk2MdaAkZXc4y2rhYUKmcJ0yC/tKH4mSE5JUu+poufhvLhmg/oPJ8bw0j14pasYJKX4e/1yAzzl9ZXz0Nh6HvIWtMVwTRidq297Pt2DytKy9d8yhhv3owk/y3EM9zoTCG8uReJmjhHUiCdfTx/rOC4ZjeT639r39iFpnzPKmHeu30Nx3ipMPgwevDluGzX7fVCuYqTDG7B3quhSw2DVv3o8uoM+qzkJg5MOIhoTdqWo5JNoMllH07qyArHzoIe3CYxbxNCiJg4293K1Snfsao+JRj/38DBQ2oII4fWHzF5KUiRY8BxFLlUbkM1T5UIcT7Z80OgvPNQ2EoNadcsvSYY88RFrmuPVPb+JEnCEqaB+oJKuUPeIPFGl29mSNYtb700JJyAlZpzJ47Ou+EYmGREwnHWIEHXJPlcTVgYqUOUbGzQRbwkt4wWJe5wHpnNoy2RgtFz7w1rRbulnHc3v60Gvkdn9Ubev0dFG7E626Dm8QAJ/ihXctVq1BZZqoXReoFVpofkKJFCB6trm8DrKvnPysn5Fmw1kJpT5jGRk6ELG71+NC41BgyjSTc+qstIkZedN8BJz60FRXblJKseWyg2GN9n89KOhrR1P5JHAtAfLhb2gMk2Dqk4DSZeAcxKUTLOZnOeHkNWFubuDM7regGbglCAN88NoZbsjUC/k8KlTcjK2d5MVwvDa9KXVpzPzcT1nSxtt5XKK28cwjUYdSZOlYro7FFsIM6eg2lBMQTL1w+ES6v5ieYKynI76aw2OMYIx+cH4VtGkx2ovYZcj9Sap5Rc9DmpnO+rIybX9fC833zjFtLWZj5LtzMgtZE2Vhsx8jnMFGVW5Kxv4gauZ3Woteazj51IzkkONGEXJ9MVncwVYpo65ZPVoFKUufV86+jWfFfPeXYWbzD8uSVz4nBipOqDVdJED0tmhMh0yiTZhUJEfd7sCs2Z/7TcZaUbLEX3aESyZ9zIf1M34IozYqnU/Fg8vt5uhDMBWROydFCL4dOh71aFW0G4Yz1hUSnE/Mzq8JuvfXRV5e14QvIBAf1OF4hMemT34mjNW+nFD0PxOHQ9WpwK7TmLrzoKOotS+QexcKFIzLJkVjE6iFn1DU59TqRKzSsS0FYX0DMvCTjHFogONx7rLJelo0nMEARCRO3q6Eo0YqvUah+lJ0HSCVhLc1Jj7HlfT1UUKLRE8radXiLGvq7K3oFB4k7CMmxpkbdNzM+qJWDARPOidV/Y6SxVIZ5kmLSa2x7rxLVrbmiVZdh6pZw5SiW+RHhy7FwnEeY6Hzf0jBWerD1SqfddYRoBBufP46kiJC23B1xNzZ9aMx4ZkDJiLsvvHKcgeipZqWetg61WHF11HVbKMGGvuhSG4LMqiEPZndD3az90VAvDZRmuuo5kxJGnXQf2/0NvjoLpSIZuhu+UfnjnnA8Yg6r9z2Sm3/RlbZ3Zx9FNOqgJrRxsuYlGGgu0hZIf2W7Pvlo3jrZ37OhNHE2u4R7KpWUF2CZdGW59b1rDuUhOn93QWRNULvmolKmsUCMVA8a4b761t1VboOGjlulrN4RQGHomv+brZKbQms45gXEFfVLDz14jIUS7cz6+ckBV3h5GWnwMecdCGYXa0HKhIkNmPyb7SphQFDfQPwXd66aMHOX20/Q7VkabEbTmhKLSrmvTJCKG/HT40f1VGD1BhX277SMPWZ5uRETgul40JinqKzQ3VOiRlt++Yu+7apsgd+/VOmKslya5uRe3LXCY3p/lNqDxvRu2AppL37N72fPJfhoROPf1jMQ7uMZmBYC9OzW6Lfh1vQC0XDsUr5V2buKTR8kVhOuoQXSXIxY9ZZ1VEt3wd8fWfchjBPFbJlj+a5ImzZCPjSImgZBS8G/EwtFds5qYYwcnwv6JdqCrQ0LLuxDCyfeXXa1xs9P3GmniCvNJgANk8Cg6zLzk/Srdu5HJ3nLX0GNfHRYrBWnhoqg9OoxNJcBn9Xmhbj9QiVWd/hwjvX4bqpYbd0moVie0XftZ65yxAYYpufYzvJl9zd4U5MFqjHZluEl0gloJZik/OLqj09UQgPq+2UCtrIQpb8L6brXgr3Rm8Vt7d31Tf67Xi5XGaxw8LOPRKALZAL7FlifzQUiT80sXhPLThY+c7772LFIshdjKLdOv5Qb2cmp4b/BNI9S/ZzLTuZ5dRzlG4LrqKEX68HfDBVzXRq4LZ8QRBX3u1mNGM1YctwKhyjQ8wdLlI05ZJuYmHOA5F0Xeqe9iL6IseZD8vO6Qlr5wLC2Ysye7ACxWC2c2JGxYfEM5GOX2gZnaSmgaYOmvG6CovwEjGAMWc+OwIYz6gAbPFFkNKQsh0Y0g0Vb6JGQBaMWIYoQEGpDwOWbxFkk0u1csTOKdbNUStvxyC9Y53lfzNbht4rx3DNew3LYqR/BGXutNjXE5I5GH8dJlY65C90Ys6w77xjWeajrcovGKHOXZGp3kpu8MBR+lMIRmy2bcQvycq+D693OKFIVL7ZX8FcyWneQ557PR5DqR3XPzYLbtKxng2Ts8xpFGgBbfBLPyWSX/04CRjM/tZkN0kZLFh1kt/IIkePDcnxNo4hgIHMdZyAJMHJxJgTXGCwvnimMT5lMIZSmjhrii2r9pesdCHXFio7peYSoDPSQ38PKgwbywmXnpjezU7VfXEMYNLHQHqFXfRfeM0H+MbIh4XVIk7JMIQL46D5fh+BG2HEd3JiJvwXHSfpP3SaSEhLCXrL6FnBzF0lzWZq7CtmMd8o+VAZpMv2+tP+Z5pplzzlzh+JObyvGW0IbkOOqYOx/rSNfUESuUUgsqo0tKSx+QgPHV1D20CUxjSEkuWvDgoUBQX4qSp611E7qL+oObQtOhl557sL8qnLNCPgNWNCsOxOIhWz2bEd1ZrQ2j2ihsKTYp17QLCl1V0q3Xpfhak9Um3TeFThQYgMv8sRCsMJ57UbLg0DmvdfUBzL0Ucolu1bV8Xiq+GDlHMoyBc+cVGIetakOObLBNeNwlt1uI7hITq7r3oQEL+bXPjwsHZsjILDC9zqYqLWgkIGXZybyXQBzMINX3+oHTcK3WgxqZioz9GNBwkJvQ/Atfv0ZehBrxppEMr715ZimsaDUG8j58TRvFVjjJS9D9GqJW6OYhZad5advlE9JGaI3rMnkeAVyujxVP/ZOVsR0JUx8Iu1BlOVPXIFlHF9LrwYxZS2rxTrPhULdfjESd0HaBqofPxjVNnnE6Ik58PiInNM8zszqzZbfObimCsdblakPX8xO+vqs+aTAYAdxj/ZzzUYTrk1yXW61HeKxcg5qv7oHSNTUYn9F5rorK9HzTU8XgLZBaJ45/52XiPbQ7PF8DJd5l0qoNyIH2ak+fXoDd9+cCe/HNRs++AiPU1lHYsoAmNzE0Vza5k81B0I/H0Oyswsxt8oiuUcDVpVPZUMno+hjEZQDkQKjSuCmomSlMCqKmBSYiypLIz6TQm6ici0aLkLrPbivcC0reo5WEQp/wYbtefLSLxblpJQiiJOj7Md7XRks6NHkTVsD9NEWuSchbuUjXe8NOQzIVtOagHXVFqVq4yXHMtWSjIslFPSwYQaFxCGQd3LNaNfYzlZADeV3ORRlKJHqt2JLQm4Drp+2g51L25U1hOMpDdErDYrlpZZCX5LpoqN0ukbkGrp2jQdGKH/05N5eSEcoLB0y8Fql76fvi+IYC8HNQmVLxw4okd7kwcXj9XylCytRuWamTgVqcOuZQ4cjgK07jRVbySMcaFepiJp8MzoA7LW5gtVy9QB+M/0an0nJPtgKKTjfK+tBMQa7fs/PrSyGxynPhzsDvttTqjZIUlGGtWolZEWzEVJhDMztknBpTIrUZHPaFUAl/53yEND/904WpaKIVAmG2oydUWlGLHuEoDCF5I7Yi7mKM0eiG91raoBiKhTC3x5KBiRgJSJraw5UPsIBrBfS8/JGV7XXzgTfOjyD0lRuZViTimzqpSdGNXstJxDOaVkannu9xvQwLWjNcc+du8tkwX6d6ZfXuuBmo7J4RHNM6VJuRQKGjtFJbPVmKMgx5SFCpcI4I/U2eGjGWu8TjAVgXVHPv7OXiwWq9FNGBE9x8H0bSGtEOA6lJfbX+EcVZ5DFOU+qETgmLzkEIpnrfMzhpWUjysb6eO59KBpmKEJTxGlav2+Nt1nJoI16KmSNS6FybYBtB7LxwivUdWmuIqjb9gHXUzBeLwpJtzIyAZAEHbJvwMLGhAt5+1p0Vc6/fLzHvpdSsdGrDoCGsXSc0VN6jg5gJXis5wG6adWF2HB0oJAEwM5KfKGvUZ3gshs4InWuz7/QhTBS9crFyIIRZDdqwvDM3ywqPlOkWVUaCKAtcBz7HXD8aBaBcvZVk+UdfzJ4TN1iiH75VqCsOhps2KA8115UfUs/FbNnQ/e2SUVMKDSU3VycfNlphdAdINTSu+9udUVm/5AxjDmzfmYS4QaRB9ORnZ8Rq999EGP5crdAxEDPXeUUA4YO3U5Eanw+0InCyeQz9bPSGWwuIOBxW6ZtZyIqxXnFgRwlHhZAOXKiNcvR5oExIOtbZyUheZArn3hVhefCIgIa+B3z2yP1AGsNuWqVj1QEwgcBjPxfk224lz/EceNKmU63GCh1pwNz8avpRix39Xi1yaVomKNG3nDn+hJ7n8aYV7FJVbQlvalF3bhzxBFbimjBrNDfITTp+lV68pNgT5H9aseSd+6HwqYfDQCiEypwTzusKczJyk7R5OllMCNKNcpCHk4LGHKNdp0PVn9NSXprzKx9au2MZgVl2dnMEjyHQlNFOmGtIzobJDgeGrjc5J6Wi553wTKTkLyLwiBcZD7eQXN0H9oHIUNIi368l6GQ7AI8LWOtJ8sIetysOrFz1TAGNuZKyXiQ7lYbOzGZIFgsFLXdpGK7UfEbK5wJJ33qF+5zcWXbGafTr54pVA1xLB/bMpA7LN32ozSBdC5W7VO18VFiMqCAhqCnk0NclT0LWlQktlQxFgs2w+HE9y5L2WiKGMF/7gZ3O1iz3o2tUOt5Dy3Ptl9qAsvChBQMhbI+Om162NVYvUOBqi5MAkidt5R3CPbKUDRsEx7imFXQhXypmtr/jJlPJfy92TDIx7Y+W4i+X0FEYWklzImV1+Dw15MpqZY9IIkYKXQsBIXW6VduWpW2l00aEh2bLNWgRckQLbdXqmagoM2pjcL5yZ2+W7Q3cbtS1XxSWpYiyBoe/X3g2SS00RGV/yKXhV7TGtQAAEcFJREFUObJu/JzYcTXCumCf32tzJsn7wMqr80+2xlLuWYLcgg47ImLsSdAGDnbCL+QkjD2+m1lUOlDnq2qN89JzEpHJ9Wg3xu5cyIO4rS/XGJ0R2oEAEubntS9ceFSxE5xuXTfk93shPXzQhfADtQKIwE2Lh/005kqsOHBx4K21VpeoJwwZuWho68M700qVr5l6sGqMU7/vFqyZK8C+EhXqPJCRDPkXMuFrudtCHEWwya/2JNN61X0aDFbIAwzXKS8gZji43IPyoJqoSyf2ZHrxIv29pABo0wa42lJPiYLeSLB/pfEbicuR8EVl3a7DjFSoniSZ/UlF/4BwSub9gByOJqHvqu8nryu3phv9jvmiNKloC7Xh6PZJ0aFgMTu7ydFs3RvdMYuFVbmZFhDKxKT/77T5SrzKGMWNiNtBT7TkiOKLomE88yhq4zP/pg9TpkLu+TpYZtD3LM16uUGS9p9duyo7sGENKmPQVdtC1L0Zwdr43Bt7kx7ofZvMtjXBK7TaSOoa8p65kWuXGwIJKDkEKwbmH7jNeI4b07rZt6eGma9nZwnaYE1Ow9CoSBpx8H0djouvDros0ZPfvnX7XzwgMTAhvQmlu5b1axy/cxD4fshdAEZiFTBgcTepHSduqb8AN3zu4T3NqIrLm4kWXm88mQGUIJAPudfMJOi6SKkODmj63k4hhmoTQute/jsb40SqXxIyqWTahhFJdhBd3A7vurdkSWsK5xA4fflOOBeC6Dnu5+DmpHa0EULLz9Kz8CeGu1sGITXnjhwYC96v1zJFpSLf38qbCof9UThf7Ki2Oe/gKX0sbrPC9rPVXLAxMefKXFYXJWZ3dbc1BzkTIQrycgBSbs7yYVjtXuxBCCsLECnC3QoIOI94gg/s4UJqiRAoC/uSL/CRf2i4xNJthpVGRl+4zl5FOq36a7IYcaFf6U5Ax3oa1mIjM3RdKrU67ChaoJYmo/DLgYsSpYxKZmSOLEsJx0jdlp+HsaD21Z1U1dGVJtpKoKHv8V4UxCmMxEcMYQKuv6DSMv9huFpCuvVaWb1SmKxiLQEdsLKfgF2iAqeFiBZ2hMZpaZwVyQxboyuey8KNcnXOAlAdxxklg45ZsDvpHIRoRBdam0r7Zpi7Rmg5GoR4LPnbM1xtqe3PSGm/il7JsKw2W8ygtNGI/pdaTs7ZzKsN1XlX2kQ1cxytYC07lIhBzGpuvfZEDfz3AnttjlaEINfEWq427L3vak0eJoKjERcqt6XW79R1nDT3xhKSTCPozibsVnz/kxq8uIP2FdeYPE7C1PKapmab2UGYGZyMw6+RP3fErN8g0tk9eAqtEcEaW9D3o8JoawBnhBLCurANP+V+dytMpv9o/3ZOejYTzvtR1ULXrfmato9zxd5IwHh/Wik+X1s1biquk5LXLL3opP2ep7iPidZ7IhowutNrzTW/jZeh2/vr/LdlgM/uz3HjeZx+v8je2sDHOjTuo9PDOUev5amebZ6HWs++QoH4XudOeBpjXsH78kxc10v4PkEKqR+TNSewConq1cEKas5H6tl7znI8bwSUsxFzj80MzLnWU3ENPJ3u/8EsYiq5uQciAmePz7OYGhP/5Fibm6LteS059hXORCW+uGqQD3iMyeTBtO3T9I3ZfKSq8tBCCPlC3H67yR8iEJ5AZlFjwkoNktmKgBN5Ck0406yUFsfI8GE1hq1TrPqU6hE/vnoieeCvLVK7GIsJKsCVL0OgXENR7y9BXt4jX2VdZkN6n0vZdQ6bVpIIhCXFpz6r+ghkk2QU7oaZmPkctcBcw1qPTn4aBPUtsaqVT+4LuXCfh278A/YiSZd63xRlC+r0hTGel5tg1nTwGjMhjRW+RWyf7fLc81q46vWZvtd+wbUfnQqduo/DfiWXVBxXBjDmzevUch3MOeiDu6kQex6gk+s9B6zMPjrCtHftF0UjwDk0wVnPvC3/4pHQPWWYIAjtMyiNyQWX9sjKbd3c4BG49oVrM3Fvy8XJoQusRid6JtnvBjk0wBtVmibrgSF8Ij82D7Edgj9gH5NQfGNfS4ojAeY/UDAMyy49jODtcImsva1p+cMNxQ0hvxkJnnXiWDqFg5uCi5VaSFYIzpwKr2j6OfhMnDM9vYvV5iiNsGY+y0ixFck3oSvvObgNcQoY7/M1Ki4rKyBbgGsM9FfZnGi6FKAPPAjVAHpsJsG4/mT++1WvU27/Pp8z+TsbsdR3LvaUpDKT8PraMa4z3Y0ZqjZXUXOihKbX4xocxhyjc2Y6JZ2+P5z/YXeQ9/R8csyAmBcoAY13HEp1ooqZjIfbXsIr5ZaaK89r/sQ90RyGM01fG66UYt2S51Y92wrtjrgTJzd8NdVwIw42h6n48lKeA0ukfaHAuZ7kV3JTzMpDgHDehUlbFsoQvaIkhMnlmlzD7ZGfjKXT0Urt1rwR3nNaoxOSmNW3xiZmbHprUc0mR69VCeOAszF82gisPqiZG1R+tK9SPjgzSNOHP6PHR8HRuOA4/ZVGCxSmNTI/9ZQZXWnIsyW44cwVlU/N7L1CF9nuy25ktBqNACyIaz5FiKtGcSw6LfSfzXlhPQ0ZaMUMpkVTLuZmYDWnG8IgGeoNH4RNF3BETWjcvKH49NfgYrzpaE9prNY6KtwYbEM3HEZGOrBu5Kb/W5pDFkcyN8RzHhqjeUE6fcz4XV1SMHgu3duuSjb5GAjviy7qCwDTRd7hwkY+O0vrE8yvOK2sdOJZ6JlAOelI11pn5anS8hJ2IPo4N1m8KoXdwXr77FLXQ1CHmni22B9kcyun1L0mjJPHmJNg6g2rpemQaCuYAwtrEKO3Tt3jnNXAIfJJbftyVwZbpjsG5dYEM9uuBMJooAQxZH2V7xDkEQa4CzeE5UnYbn47Q2SNdsIpvDyKkX6qLSyFbzXPbNdRqeayXIPUa+vCZSBUlWKjFWWuCCCoHBEQCBuKrWpwAKwEz6aImE1UnCfA2WNEq6B/GDWJYOS6h0g+pjBTjigrlRFrtmG1UmFBn09fWwi4TaE4IYbqm7BXSTfcSkEHWzXXYR8fIJydBmzDRqgygQ9tzodC1yqikDyQAEVidEPXtA202Ahmt7rZW6nYcx/n3tg8QDqrtkYTSJSYXh+iCyZDClkTpKA8jDOxo3wUCkg9JCK0AXe+iKmnwDVgQ6YFqxZ3wvmRvYdK4JkbQ/0Ewe5GZ6ddU0vyQRawEkyJVof//VwTHVHCC0BdruBJhngPRjku5YOIc8h08w8U57Fa428pQbphAJpFdkJNM9I8n2PAt3pOVyzSZ2dePze3e1125iChYNkO0K0zV54SCPMlG9feiPAcFJrpRU9u29pqOqhYyq02dMlure8RM/+mG+oocsIM1ANsXJOSTSOmOd9TaKmQLmbuYuZdzDXk83LOqnBxjxZ/AuO9EbgEbtYDKcmdtY15Dkv23PD82orymGtia8TdSGQmSZXKOjV/uZlVmi3nS6tV8+yCMa5JzRb337o9t3kfN9Phz2453ejzeoIRM8r2hWqXQdmvLFWXUizvF1zKO6qkuhxKP+NEZh4dGtmAUpINo0pb7thakLKStqIrFs44sZEd1QgtggQA7hvJ67/ur8DjDtELu+LECrOyR4yCoW4espvYQzxZq9MC8l4kbeBGMCpmIqE1wn/mVKoH59EQf2ci+3sMt57xpA1WTP5MHqvxnJ0qbL86RA5TwAOhhLAjKt2XROUMZbL/BoEikRe5nsCJWFsKYQb+jjjVVV1wWmgkQAPkXqXe8IoqpREaE5VGHAbB4wsFi4cSDFJ3pe3rpPGWt/UE5aOE65CSpf/hMVSi2DmQg1agd1dhD3tqqXWJNdfBz3LEU0H6dLm70c0SIsnMarXAay+7r8dy+jot9VGVkI2gaw7WwVPjqUTqv9mkya6Bk9Hqv9F3JVYnOzOy1L10RypD9DGjVzLv0wj8XE8lY5JKpjNYGTk5EnlW2zOSRrCFC4rxxoonQRz9JLp0uLS0tRNToElMsQOWE03Qr9s6knF2D8PyLR/mA8RYk5ADVrBPwdmT3638ADxYXyBrDR0HsHNXu3+wdVkTnsuWuuLKh0jBZIUiYiyiUQKjFdWmzhPOqAwFRjkIN6QVGpdsAK/Rf7Ooq9AJN019+h5ZMuKrn91qa5CWCAAXkJNj6VwPPF59zv+f3I6JtPo7FqEw1wjI8XxOSx7Ebkuci7RYiAXYMpr8vPYLlKINogA2zgk8mGeQHZXo8VRK90x02lqHndugjEgAjbY603HnRqwTV5alvvgahls41u+WB7EZsufne4WGcar9sNXwV3LbxmwJS5YCVnElXH5B5cxESSojEb1jTaCj0Oj6cRe2oQZdbRrOQvknGV3ClM2JhkMnhOla7LbEK9kVimtNpRGoQjMrF/u6KW6ABNBM5ZXvP1n5sZmIQnhAbnThjzzZWwJP8x26fmtguKeDyKk+N6TAaY30iKPdHyc8laCdFjwqVt6jxz5dFBFXaauQ6rptBTqThQCohRs3JPtaUvs7RyAwLiPBF+SnPSc8HyvCOWaIsoi2WmO6DexiJQVPN7M3Xglo6Mrt64AhTLPyIWViq10IkgqPZ7UY1YbkJBrhxXgCVf/GQDzDesqdoVILVnQaFQm1lanTd0jsEiWsyHJHNN+e9GOdCq9OdCv+Y5CtJPonZ0XUxLDxahTGvKTd4X4QoSBB3otGneSxUEhACp3qwK9VGz4/tz2FRIo3m3J0BtBkUGtxNPRIwneAx99Vdlh/BqHU7Mpoa8KwsWzWaMCy79zZ5w5nWXCSav2gdabmSC9Pl5tHL0ZIULkZO8SFyxtkWHJbyLK0sRrF8NzMsVA7N3IxbNSMTJcW73111ak31dzkJazulEVLlahKw0efaYJM7MuhYgrWxvaBRgilSLsQqAW+8wnAk9v7mReKsJQLyU2RJISdWq1MW2qN5CYKNScSUdnjU61FW9IpJ0joCL9pwbBfRZdQriWjBUIY0VzBHh3UdveS0GeYc/OQAVo0ZmiF102BRcg12jE6TTrj/Yyd2pzZfElHHGj4ir1F91PAvh4aAyM2vB6i81NoWINGzp3h1LYxoQrSOgUvtQ6xDugM0oTQIMP6zEPybQPYV9Xn0Dsooq9cqnbrY1Uti5DaGgo7s3t7QC4QjR5k7Op754rjReXVjQ5kCXulI+IWOl2xEOsJieI4Mit0Wm5JW/22NAmSXzxuHn4N1HLOtCyNTyvOkBGFziFE++1THCF4rk5FvAU3tWAurUPKn6t/+Zc68t5JXeQ7eP8Wy9pIN7Z8pDWnM1hn8A0xLJgIrbqqIkqwT857blQT1nIfefBN9dOQdWrXKxt5EVaSgygnqF/r9bqSmzVuVo7/7hnVGtAyx9jMQFRfj7jnlHDuyy+fh0V5LY846YlITtAcGaNV5Eio0NaQAK51cKPzWSNupQRc3Nmmj+u74sDLflZEZCY0yTiwSRPvrGfnMIgincb/GsWpnD2G1ClKsyywQtqd3dobWakJsYSIEX24UCOR86g2DMc6S5526pQ4rucRB1g3Kxkm2R+vuJc4Xs7PXn7wt+Mp/vsVx1NaJGK1Gd5xIWLlta+44sjMC9c64sqNAysRwIV6b+cV5zo3gLg6H+Oi73S84CV+HIHMzi6MiMjMXTYtMlacWS3lF2Uoc2esVWdSragSasfVo6sETzzwjBpzXS4z45aVGiRUgX1dcRxPScVBi87cgmxkdEVgL8LQlVm001h6cR7xiKUz0pFQtWVB7LZKrSSZaYoAzngy5xC2/uXqPWLFSidLrZZWICKansmo7FPgwNG7L2NnzTDTjM915i17szZvaS26nZHd8T4TUL1MtEughJdrq6AuNZ5ulr+xRQ8Ckdrc2gNd1t5fWdUHM6LDX0ITa5V07CsijuzMzVhYWTkhZyHKsZkVYqSVLGWTuXa8RoJr+XCmMo6VBvDAy41IjTiw44Ednxfwj4uYLoARZozVY424YmXxU52r0pIz3ctctXnLyjexrXyWliSR21SWiJ07V5yqjr1yR6fOZ0YdwrLjwl5nzXZsXLHiwgOsezrWmTs3drB1ZYLAEu0+rliRidx5xbHW82eff/9v//9C1gNRQJVi3wAAAABJRU5ErkJggg=="},{"background-color":"linear-gradient(to bottom, #ffffff 0%, #ffffff 100%)", "background-pattern":"/usr/share/com.github.philip-scott.spice-up/assets/patterns/bright-squares.png" , "items": [ {"x": -201,"y": 50,"w": 878,"h": 320,"type":"text","text": "Page Title ","font": "raleway","color": "#861002","font-size": 28, "font-style":"regular", "justification": 3 }, {"x": -202,"y": 314,"w": 1951,"h": 728,"type":"text","text": "Lorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim venia, quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo consequat ","font": "open sans","color": "#666666","font-size": 16, "font-style":"light", "justification": 3 }, {"x": 1447,"y": -385,"w": 176,"h": 585,
            "type": "color",
            "background_color": "linear-gradient(to bottom, #ef5b5b 0%, #861002 100%)"
         }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOy9eXBly33f9+lzzt1xse87ZsXsAwz1uIiiVsZmpEhRtLkYRwwjV0UhTanksqWYSaTICZPYZecPSxGdlC3ZScWuskuuSKJkkRJXke/NhsFggJnBYDDYgYsdd9/P6fxxb1/0PTiYt8x7j+8N0VXAvfecXn6/b//Or3/9O7/uFl/84hf/x7Nnz37WsqwAYBiGgTs5jmMbhiFkJQmVp1wuI4TAMAwcx0EIgZQS0zSRUtZ+SymlqCQDQEopq2Wk+u04DoZhqDISQAghqiQIwKn+llJKQ9VdbVdKKYVlWVTro1pFjQ53qtIgtDxGtU1s23ZU+6ZpGqo+x3HKKo/jOBp5SI3OEwxfEgz3/v6vNchE4ighbzD5zo+Wm37113PvdwwdxynNzs7+rnXu3LnPXr58uR2gUCjUGFKAOY6D3+/3BMO27VqlqpyUEkVAleHaPfXdcRx8Pl9NGE3TrOXX63Ecp/bd5/PV2ioWi7Xvekeodg3DwLbtOnpUXr2c+g1QKpXqfqvv5XK5Vk8wGKzVp/Lr9J9g+HJh+B3LoiAdzzbfSAo3NFijo6NRnZ73K4a2bX/GMk3T7yZOJSVoOmN6hTqz+nelnfR0XH43iG7wVB71W2dEv+c4Th1YXvS66TyONvdDpOjT63B/P27kOMHw/YuhIyXOCygL3Tp7v2NoWZbfMgzDLJVKCCHw+Xy1zH6/v1ZIaTU38ZZleRKsRighBMVisdawZVm1vMpEBCgWizVgVbtCiJrgmqZJOp2uta+0oxoZVNJHS0WHPrJKKQmFQrX7mUym1gGmadaNNnoHHfdwqeuKxxMMXy4MHcehOkN5S8m27TpF/H7GUEqJJaWUbtMVeF2NrF/XK3cz49aI+jWV3NrQzYii77iR0g2ae4Rwt62Sbqa6O1Qv65Xco/QJhi8fho50XsyycP9+H2MIYOkVKjB1ZgzDqGNGN2fcv49rXGfeTcTzTCovxnXi3UzrjhlF23HtqWs6z/p9r051m21unk8wfLkwrExD3rploRTNy4AhgCWEcAKBQM0UUZkLhULN9CmVSke0shD1TiM1lXEcp2ZiAYTD4VqduVyull+1BdRML51wwzDI5/O1OsPhcA10HUBd2QWDwVo9ytxy16/qdHeI3nFSyqoJWu8Q0j3FymQFCAaDtbInGL48GCoe3moSQtT5gN7PGJqmiaUT5jZbdaaP+zwur0q6VtWBcCf3Nd1ErL6+8TTL3COol6Z10+HWpCqpTlB5vRxKx/F5gmElvUwYvvA0xKP+9zOGtWmIIvw4hnUCFTNe99yNuBnzIk4XUj3pJrFywBzXlpf55s6n53XTrneaTstxQCtTT6fzBMOXC0PHedFpyFGl+37G0NIDQnSTRidUf/+sm6bKY6wDLqWkUCgcAcf93l7lVX+K8XA4XLume/WVaSSlrPPeqzqBOvNSZ173DCtzVPGr6FP1e/GiP2w6X27tfYLhy4ahg3yBaUi5XK69oXi/YyilNCw4ahq503Fax20+uc0YKesdNwoEvZzXffVddar+2kinw61BtejFOjC9aH4en+7RRm/L3THq/gmGLx+GL+rg1Ol4v2MI1WmIeyTRidJ/H1exVyNeppCqX/fIquu6SabAcHt0nzd30ztap0MFGnk9SPr343jx4t/dObrj6gTDlwdD+Tb4LF4WDKWU0pJSOmouq1emzCGgjkl13+0w0kcuvaxu0qjOkVLWhdwqk0yVdTMiRL2TR6dVjZzKY6zuKVNND7rR52bqu96Rbu0sxGEwj/IMq/Z1L7e+nuIEw5cHQ9uRvEhQlkS+NBhKKYV1nDZzmzvqmiLmOG3trkP/7h7d9OvuMvp1fYTQ35V71eOmQxcSL57cD48XXfqDdhyvXukEw/c3hi9qWTjHYPR+xBDAcs+dvMwYdyW6wOnEuOtxM6U6ya1N3Xl1UL0YOM6kOg4Et3f5uPJeHeUO5HmeuXiC4cuF4YuuDdF5hvc3hkIILMBQnladIN1bbllWDUzdc657U3UPs+5xVd+lrPfieq2u0xkRomJ6qVc7KuAEqF3XGXQDoptbeicpzzNQV4cy/4QQNQ+w4zg0NzfXRqFUKlUr615P4W7rBMOXAUMH+QLTELef4v2MISAtRbz+WbvrGql0raMnd3n3HEhpcrf5p4RYn6e561U0FLYXWPrma9X6JSDxt/bQ86EP4w8F6sxnt+nm/vTS1Dq/+m+Vz619448n2JqZRapyUsNMQLDrFCMfvcbNL/zPXP61f0BTs0kpsY8RjCLMSv2ZuQkef22GVz7z6XcFQ/27ez2C3sa7heFxo+t7RQ4dKbFfcBrysmAohBCGl/mjM6N/P87sOa5BnenjTKPn1amXST+7ze1/9n+Rjm2Q2dwgu7nB6h//Pn/6X36K9EHmWLNT7wydz+fxpIRJCFHn7FHJcRxK6QTpjfXK3/oSE//wt9mZXSCzuU4mtkF2/wCQ5Ha2kE6Frskv/CqPv3K3Vk9xb4O1W5PvGoZuHHRHnzvvu4Ghns9dVqf/uyWHlaAs5y3/SXnI48uAoQVI3QwCamsKVNJNFP1VnJeZB4ehxW5TR0Wbuedd+jRIbewhRCVoRNFWLtsEB0e59plfqwsuevo7v87dL/4+P/T5z9XaUF59RZviRY92U/UrIPQl27pXuVAo1HWYGoW6P/Rxuj/0cYQQFPNxVv7o/2P0F3+FtsForf5CschH/vEXAYdcLkfZtikW8nVzZqF14DuNof6WRMdQD9x6NzHU1y/oZvl7SQ5fZBpi2/U8vp8xBBxLH0Xc5owOpJ5P3VcEK4ZU8jKt3PM3lXRz0N1+XXv6f00zjvzk32Dmc/8bZedvQy7Oypf/mNi9+wgzyMDHf4rTP/KxwzZKeZa//IesfPsmZkM7Z37uF/FnV9jYKHH1P/1Ehc5ckqd/+P8Suz+NEW5m+Cd+nr4bV49goISqRkt1JlLXWU6WiX/0D7n4K7/J9h//Hqt3pzGX/yn7r32J7/v8b1XyurAoJ3eZ/8N/zfbjOXzNXZz56U/SefHM24OhR//q+dxWh9vCcMclqHy6aa/u6zsv6e09D8P3mhy++BL1o2843q8YCiGE4TZf3OaZ+q48xzrj7jz6p9vU8TJ/dM3uZUqpcm7GdHrsYh5MH4aAh7/3v5DJB7j4S5/j2n/xSZ7+83/A/X/35xVAywXu/tZ/zYM//CpDP/ELDP/gh3j4u7/FzL/99+zMzVfASu/w5U//LAcHBtf+m7/D6E99gidf/E3u/5s/OoJJPT8VP4XQ7gFIu8j6N/+SUsGh96//PJ2jp+n9+C8w9pnPEAj7j9RZ2FnkK7/0SbK0cv2zf5ezH/8BJr/wOR7/h7+qKaIXxVAXFoWhOzBHv+cloDrdesyAUjBK+I6j93kyod9z53+35VBFcL7lv5cIQymltAChzCJdkx3nQdU1ozJ7lLZWDejLXXWi3UIJFc+rbjbrr7D8fn8dGJWBWBwuxXVKTP/rf8nAX/txAn4/Y7/xj2vtlctlXvmNv8effv7/5OJP/QgHt77E0kyan/p3/5ZAsGK6DX7sR/nqL/0nWL1XSSQSzP0fv43v2k9y45f/q0r9A4P88O/8C/70kz/L0A//IO19rTW69V2nfKas4+eQfh8CgWlZNHYOEIpGCHX1036mYinkqhg7UoLj8PB3fpuun/zb3PjFn6rgMDTMj/zuab70Nz/NwEe+RKQx+EIY6iaovpxZNzuVuS6EqDNf1WjsFjK1h6VhGCQSidooGQgE6vJ4yVUdhj4f7zU5/I9+7w+wSyUqvge9rKz9FkJZDIcYqjyBxuaXCUNhwdFdkVQFiqnjnDP6d10L6V5mdc/dabpAe71DPtIGkH50i7/83C8hqIzm2fUlzK5L/Nj/8DcrnVTIsPHtr7H/bAkRCNPQ3Ux5L44jJRt/9XWGfuIXCIZ8NeEQgTCDP/JRYnsgKLP+jVcZ+ZWfJbW2UtfB3ZeGWP3OBG0/92N1PLg1uttkrd1TPB4zsgBIJ8fK1yf4wE//vUr7UtasiY7hBtbuPmH0R6+/GIb1I4Vn3+l51W8vy0Rh6ObX6+H0ossLw/eaHHZev1Hj061w3bzpc363f+RlwBDA0ivUC3qZsyqfO4DlODPILZy6910XxOdFpdXyAcH+M1z59C+jNLvV0Ezb2XOYloGT3+frn/kUzR/8SYY/9mM4xSw7d75WWyZs5wr4BhqPPhhCVN56SptStsDSH/5LtpsPN0oxhIGUUdo6okdogqqzyqyQ5Maw1jGHgNRhqAGFoEwxk+PJv/o9/EGrfku2hiEiTf4XxtD9vQ5fTaB0PvS+c5uretlDVryXXbvrPoKhZnLrZd9rcvi9iiFQ/zbE/V5aFdbNFXcQi9dopf9WppfuQNEJVd5aVZ/7rAdFU6lcxmxopeXytbrNTm3bxrZttr/9JxSaLnPtlz6FqNbT3NvEvT/4KsVCkZYrV5j66l8y9slP1ExHgNzWDtLoJBBqpOPSCM3/8ae5/OM/UFe/m3egRoOUEmmXQYAh6jsLp14QhRAY5uH27cpclVKCiNBxsY+R//xXOPXBC3Ud7RXY85Yw1N6AuDFU9emmuz5aqgAhIcSRNQjqMxAIHOl3t8zo9NdhqMnOe1oOv0cxFKJ6oIl+0ZXhiJaE+ogzr4bcmvY4TaV3lG5OuTWnlPKI89DdZrC1k/TCY4qZ6rr/Yo65f/MH2KKMdCS9f/2TWFu3uP3P/oB8Ko1TzLPypf+Hp1+7Va0LLv6tX+HxF7/A3spm9ZrDzrf+PX/xdz6PpJ4+3aSrwejSykKjUwiBMA1SywsUEvvkD+II06C4v0khmcIulLnyy7/K/X/yW6R24pU2nDLrf/LP+cv//n/VansBDMXRqZNbQNx1uEdeVUZ/kPQ2dGedV7vHY+g9cr/n5PB7FEOoRnDqJpIbBPccSNc6XuaNDoKu3Z7HiLteN9EAmD6sYOBIHpWv8eqPMvqxr/Hnv/gzNA8PYpfKnPn5T9N76zVi00sM3jjND/3e/83kP/kCf/rzv4+/uZ2Bj/8Ml372E2wlKm03XvkhPvrraV77u5/G19aDzCUg0s0r/+1vIpCH0ZpucJFYofBRoRQCKxTCrGJ4+qf/Bn/xG59n7c/+BRf+1t/n4sdfoSn8v/MnP//jXP7c/8Sln/wZXskU+Pov/wLB7gHKyV18nWf58H/3WwjxNmCo9Y8Xhu5PrzNE9Ha85MVrNHOPep4YSu8l9Oree0YO+d7EEBDiW9/6VvLcuXNRPYMu9LpWg/pt2pSXVYijJz6ppI5FcwOr59FNQ+UZdjOqvMFAXfCM8hirekqpOKV8Gaupsd7B5dg4ZQfT76sDf/offZZ8x49w41M/fQgikvzuNiIYxRcJHQHQDa4uEG8HhtIpk96MYTU044+E33UMVTv6GSLuwD0vYdfp0fl1O/HeDQzd7Z5g+GIYPnnyJGUoJtzazItg9dtNsHt+pDOiTK/anN0wPE0f9/tld/vK3NJNLnebUkqshibCHe1HBCM1+x3+/DOfZX9pHdt2cEoFdl79U5587SFnP/Fj9bwJg1BnD4FopFa/Lki6GajafjsxFIZFqLMHfyT8XcHQPYrpwqX37XGjoJ70et5NDPXrJxi+OIZQ2YPTkyk9ow6Ul0nmRZRbi6n0PGK86j+uzue16+YDIHrho3zgF+Pc+s3PkkukEaZJpP8MH/un/4qWnuY6B5WiU8dGp9tLCL8XMHyesLnzKTpPMHw5MARtd283EFCvxZRG1c8v0N8/K8+qlNLT06vMG9WO7klWuwApbV+zErR6dI2sr1lIpVKe2lQHTn1v/fAn+Gsf/YlaHmWaFovFuuXb+tsKZXYKUf+O3e1R1zvjZcYQ6s1dhaGU8gTDlxhD8NiDU2/EyzHkpTGP02bqntuc07WarjmP03Q6LXqoqupUfY6o8+OlwfU63Z5przrc9/XfOi8nGJ5g+LJjaBxnkrgLq0aPA0DP55XfzaRXWfc9Pal8eoe46z+OUZ1md343YO5OdgPmvndc+3o6wfAEQy++9fzvdQylrGzYWyuonzSta1Blrkgp63bR0ePJ9eAQnQgFqtsc00+Y1hnVA1GUeSZE/Zb22Wy2rl1lXumbr6qTsnWtqo8CbsD1JcA6oLpJpjzehmHUYaV7kk8wPMHwZcQQKmedemoiHVA139ELujvDbT551efW7m5A9I70Asxdt06X6kgv081LWx7Hh1vbqnmoDqy7k73qPcHwBMOXCUPDMCpL1N0AqN/ua6pinfHjCNXNK3Vdn+fpSQHhZb69Xv2qnDvqTV33ak9Pev16ctOv53M7inTMTjA8wfBlxdASQgilrUKhwwCkfD5/xLsrhKjbmUctf4ZDj65uegF1y2x1L7NyKAF1JpPSyoZh1M7mVNdVPZHIYfyDvhOUMrEMw9CPXavxJUTlBG2VdIeXfq6Dot/dCTr4elldQE4wPMHwZcTQMAwMXaO4idJ/642ovF4aTzehVNK1l55fMaeX1Zlya+jj6nXn0csd52l2l9M/9bZVOTcOKrl5OMHwBMOXFUMDKquhvUA4LqkKjzNb3ug1vUP0TvTK777nZSZ5Ja9IO3eHuc1EL7C8TDcvHk4wPMHQK73fMYSqg1Mxo7STe4chXSPpy2x1AN2BK4qA42LyldkmpazbQUjF5Kt2VRk9OESZiFAfw69i9d206SdK60Ev5XK5VtYdJCPl0ddj6rppmrXlzFIeLlU+wfAEw5cVQ6gEZQmonzepjMdpNC/Tya0NVdI9y+77OoHua3pSpqJiyq2dde3qRYvecXr97nmgm24verxoULSdYFifTjB8yTAEjqDifnXkTl6guhtSxHs1/EbMJLd5Vi7bnmae6kBVRgHg9V3P50XH8zpQ19JuIfFK7zSGlJKsbO55tp2Ob5PMFY9gqGOkpzeLoRrZVNk3g6Fe5ruN4VuRQ3XtuymHepl3C0MpJQYg1G5T5XIZ27YplUoEAgF8Pl9tE1AlJKqgbdtYllX7KxQKlMvl2k5CbpNKMa7q1xkwTRPTNGubidq2fQTQe5MPsHy+uqASISpe5UKhQC6Xq9Pcfr8fy7IwTROfz4dlWQSDwVrdXlpfB0YfRZT3fGVpnlL1HAl1Taf5XcUwn2J7P+mJYXIvxn46dwRDv9+P74UxDPDk6RMcp8zi0vKbxlDP82YxXF9ZIl/+7srhsRhmU8zNLxyDocHa+sbbJocvguFblUOo7sHp1q5uzam+e0Wc6fd000ifG7k1rF7O3YYXcDV6pITqtcTuBvPLm5RLJYbOjtLR3MDszATZAnT0DNLZ5Ofh7DyOdBg+e5mokWT6aQxLSAx/CNPOkyuW6Bo4TV/H4TmSx2noQ4wEc7NTpNMlbMch2tbN2eEeHs9MUyhLfMEGLpwdZGk5xvnzZ5B2kWdLawz0tHDvwSw+y4eNQYPfIJMv0NTey7lTA4g3hKHD7PQk2TIEzCIYHUjHZvbhNEVHIKwgV69crNEpywWmpmdwEISibVy5cIaVZ7MksgXK0seVS6NHBNTdFwBPH0+TK0kw/Fy7dgnDgPjWGnfvT5HNlzh3ZhikfF0MS9kkUw/nkNKmf2SUlpDNvelZLNNCCouIX5AtFGlo6eLcSD+xlWdsxzNIYXFl9DT3Ju/Se5Di/LnzRIJHnZLHyWE2scuj+WVMw+DM6GUyuyusbh4gbZtTFy7THDK4f38S0xeiXCoxMnqZRp/Ng5lZDNOguaOXkf5OnjycJl+GQEMLl8+fYm9rlaW1HYRh0RY1mHq0jCMFZ4Z7eTg9TdF2aGjpoj1kM3H/PiUbeptMMlYrXc1hsgcbxJ1GgqU9VrfjFAoO4x8Yx2++ETmsf070V8Duvny7nmXD/ZC6Cz/PVPN64PVGveZJ+ncvc87N2OFvLZ8sM/NkhRsfuMGNG9eZe/QQhGBxbZ3L18fo72nnwYMZLly5xvjYGHMPH1AupCn5mxgbH6d4sErnqUuMj11nY+HpEdC8eANIJeNIYGVtnTOXrnB9bIzd1QUKhSy76RJXr13j8oWzGNImmawcXiudMvFkEiFt4jmHa9ev0+7PU450MTY2TmprFf3Qq+dhmIg9Ix/oZHxsjJ7mKLZ02FqZw2zu58aNGwy0WjxZ2kKRPjN1n8HzVxgfG0ekYsQSBfZ312nsPsXVS+cxtG49TonjlIjtp7h2fYyxa5cwgHj8gJbOHnr7+zl3egik9+jorssXjnJ9bIyx61dZXHoGssxBzubq1au0+XM1TNLbaxQLKZY209wYH+dMTwNP1hL09fdy8eIlIkFfXb3Pl0PJ/Zk5xsZvMD4+TmNIMLe0zfj4GDduXOPhgymkdNiMpxkbH+fG9UsszD8lsbuOv6WH62PjDPd1sbU0Bw29jI+PI5Ob7GdyPH66zviNcW6MX6O3t5eegUFOD/ez/OQhjT2nqrysEGjqoLe/nwvnTlHOZcjmK6Hb5UKGTK5ALrNH3mzkxvhV/Obry6Gbb69pxtv9LINmWSgzDI4uZ9WX4qoY8ufN0dzmnfrUg1vcR6Sp8vqmqfUeae09sVPAiDRgGgYFBwJSUiiV6OjsJOSvCFI8fcDi/ByGYeALhCmWbBrCFW9xMBimIezHcUoYolwzyxT9utbVTTFZVVjhhigdzU1I6dDVGCQnwlw61cPU5CQNLZ2MDnfpx75VMPT5aGtrJeD34/cHaW6MYBgGpiGxncONe5+H4eZWjLah70NKSXN7C2YqRzKdovP8RUzTpLWjh7XHMWRDxbxN2TZt0TACSV9nG6s7CQwzQHNjqE6Q1BsBx3GIRCL1prFl8YEr57l96zV8oSYunT9d7Q+7+nno8Hs9DHc3VljbieOzBMlMnmhDhO6uLhobG/EHQjQ3VYKc/D6DUj7JQSrFgwcPkE6ZxrYBbMvE5/fht4w3Lod2gbJlYZeK2ICd38WINFdoM/2EhMAwTdrb2rBME8cfwDAFLd2nSC3Oc/f2Ov2nR4nHd0nIEveTm5RsEye7hxFtxRCHbygcx6FUKnGQTiBLa6R2AF8Yn2Xh8/vIZrMUSyWKsrL+w7EdECAdg86Oljcuh1UebdsmGo3WrIpMJvOOPcu2bQvLbY7oAqru6a9PvB5+t7bSmfIaKb3KuMu7TfC6+2YImUlRdiQ4ZXJILBeQbY1tnBm9RNhvksvlyOwuInAFmXjw/ly6qNSfTcZJFUqELdjLOQxYAl9nH21d/dyfuE2mv4tCueJgzKXiZLLl+s5AIqVTxfUYHj0wbGlpZyW2RX9jP7tbu0gaaG9pY2tji65zA+xtrRNu74R85dyTFp+PnWSOzsYgq1t7dI6eYjtO3da/Os/eOEgaW7sYG2viydQdDvLDCj0cu/7M0NfDcH55hQ995AcoZeNs3HmE4+gOv8o0U5X1h1tobdzj8uXLtTYmt+awbYk0HbZ3tuns6Hx9OTT9kMtStB0ClokRaMZJLSIBu5ilIAyEq2zFHhEMnRll0LG5eesO5we6MGQzo0Od1UwlStMLOPJcxfFnmjjligO8o6UNp3GAkZ6WSr1OEbt6zwoEyFc3ld7e2oXO9qocer9Z8ZRD1xThEMN6WXo7n2XDMDA/9alPfb6trc0P1B05f9zcSH9v+7z5tZ50a8I9L1LX9frVd30Otru1xkZsi1gsRlkEGe5tYebxLBsbW5y7eImAz6RcLtPa0oYQgs72Fh7OzLC5uUWmYNMUCWIbAZoaQhTyeaItbRg45PN5mptb6k5hUgApvhSdhUKepuZW9nY3yaczrK2v03fqPGGzzNT9KWKbmzS0dNPb3YmTTbCwvEY8W6C9vYXW5kaKNrQ2NVLMZ/GFmwj5TErFAtGWygj1ehgGIs3k9tZYWYth+8K0NzXR3d9PfGuJ5dV18jLEpbODlAo5zGCUgb4elp8+Ym09RqStn/6OZkrFPA3NrVjG4eilhzDrKxeFEDjlEg8m77G6voEINjHQ3U65VKS1rYNCYo/1nThtbW0I5OtiGLAks3MLJLNFOtpa6WxvIV+StDRFKeQyWKFGQj6TcqlES2cvIZFn9ukiW5tbRJpaaI0EmZ2bJxwJ8OjxEoMDPW9ADgXtLVEePZplc3OTSFMbnS1BHs0+ZXNrl8vXrxPwmeQLJdrb2kBK8sUSRjHL9OMnbMZiDJ4epae3j/jmEksra2zvHtDe2U1rxOLh7BybsW1au3rIH2yyk8hxbnSUzeWnrKxvsHuQoqOzk2Jij9WtfXoGhthZmSe2vQOWj5a2DgKmgxmIEvKZb0gOdZlQh1pD/aHHb/ezvL+/XxTf+MY3kufPn4+6K9Tjw9VZBsrc0c0gVc6LmddL7jmRTrA+okL9yj63qaZo03f+0evVj3LTpz/6uQnFYrHWhr7cWKdBmeu3777GB7/v+xGCYx/wEwyfj6HjHJ4A/mYxzO5tkDBa6G4OnmD4FjF8s3L45MmTlKU0l86cfk0HQQdVAeRlgrqvHceEO+l16zSoDnOXddPjTu77xzmC1OdxNOv0SCnp6uyu5vX2/p9g+PoY6tffLIah1h5CWr4TDN95OZRS4nmKutvZ4WbCTbBXI25i3Z2i5lpuhrzqdgPqBYqbB6+yOm/Hge6m012XlJKB/iFUNv1d+QmGbxxDLz5OMHzvYgiVtyFCVaTHveubguox8PobDeWh1Zlxa2GvOHMpD3f7EeLwWDc3WDpzqqzjOHWnQis6DcOo201Ip0dfF+COs1ff/X6/p3mpg6XmgbZt1+pxt3uC4QmGLyOGQlTO3ZM6GDpQKqN+zw2Cntx53MltxnnV7wbYqw13Pfs7mxS11bdeUW56+eeNPnrSO1S15/Yme40MAPH4Ps47gaFdYGN7t/6aPiqVs8R2428aQy/e3wkMs8k94tW3AXoZLwzf63KYSewQz9YrGJX2dmKU+e7L4duFoZQSQ2hX9Up1MJWJozfsJkgXQD3P8zpGZ8Zthuka00283p4Qgu3YCgUHnj55SEkebVNKyaPHj68Ya8wAACAASURBVI606aY5vbfG4uZBHd/HAXqcOah+z80/qWs3thl7WzCUdp7V2PaxGMpSitXNvTeNobSLPJp7eoQOnQZ3eS8MvWRHL58+2GQ/k3dhWGZLU4Dvphw+mHlwBEP9t8Iud7DB0tZBHQbpg20OMkVWn84QL9Q7GHc2VsjbbxzDzc3NN4yhmwf9853CUAhRmYYo00R/DaN7dPWKdc+tCprSTSAhjh7Zpr7r73JVsIfuXdbzq7bU9Z2NFbb2k/jDlcAgp5xnZnqGkiMo5Ar0OQ4N0UZMIdiMrZDYj5MtlukZPEVvRwvNLU34fD4eTk2QzpfxhaLcuHaJva01lta28IeinB1so8kOkkvusX2QIplMYQYauHBuBFnK83h+gWw6hRVq4uq1y/iMw2Ckg50Nltd3aO7o5vzpoQqGPj8trc3kUwfcvHWL0dErjJ4/cwTDYi7Fw9mnlMs2vUOn6WqN8nh6inS+RN/wGfo6W9leX2J1a5/GaKi2FkDHcG1xju2DDI0RATQjhGDl2Syx3TiRpk7OjvTVH8knJQtPH7OfzNLZP0JvW4SGSBinmGXrIE9vdxt2IU1sP0tXa4RHj+dwpKSrfwRfOcX2QZJUMkXf0Bky+zEyBZsLl6/RELRYXZhjcy9BtKWTc6cGKJeKzD95RDpfxqJI01C972Btboqbs1tcvXSRgd4Olp89IZktMnDqPG0RwbPFVdKZLL5QI00Bh+39BG3dg/S1R1lZWSKVzlN24NKVq/gMyd7mKiuxXYQZ5MLoGUQpxeJ2kkQiwenzF2ltPDzpLRIJUyxkWV5aZP8ghS3h/IVLNDWEiO/GWFzdRFgBzgy04TNAIJl7PEM6X8aUeRrDAwTCDQQsgVMu8nBmBkdY5LMFBgyDjdUlegaHkI7D9uY6XX1DbMeW2dncIV8s09k/TG9zkNdu3eTc2YtcvnIRA1k3DYH6qYT+qSsHfb3H2/0sAxW16TY5dQK8zFW3dtSdNV7a87h61Xd3Xi+t190/zNjYGFZ2m+1smZnJCfrPXebatSuk9veQwM72BraEmQf36Bo5z/Xr13g68wBbwubmBjK/w1bW5OrVq5w/PUQpe8DjpV2uj41x9dJ5yrk4u4ksmcQGmxnB2NgYYTvOTqrA1NQDTo1e5vq1i5TKTk1RCCEo5eI8XT3g+vVrhMtxlreTVcIhFlunoaWDnr4uLo6ewRBHMZyfnab37GWuj43R2drI/Mw9Qh2DXL92lbmH0xTS+zyLVUKf2yM+svlSHYaZ3RXWEzA2dp0gDraE/Y1nHJTDXL8+Rtje51nsoNauEIKNhceUgm3cuHGDtblp8sUSsa0tnGKW7d2DSv3lPJs7e6w+naZ5YJSxsXH6OlvJJjc5KPq5du06Tx+8SsfQKOPXLjBzf4r99WcclEOMj48TKu0xv3HA+rPHmE19jI2N4eRS6IOglJLegV66B4YZHuhh6fEDAu1DjI1d49GDSRy7wKPFDa5du0YgH2OrEGR8/AYbC09wcJh8NMeV69e5fvksd+7co5Q5YG4tztjYGEOdQabnlpHlDA/mK6HZTZFAXdux2Do4NpOP5rh09RpXR0d4+PgJpWycx4s7jI+Pc2n0LOVcgv1UnrX5R5hNfYyPj2Nn0yDgYCdGtuQwMzlBz+mLXL9+lfT+fkVBxDawnYqc7GxuIIGH0/fpHjnPtWtXWX42S7CxlZ6+Li5fOo8pjp/2eF1XfKh77+SzbLgfTK/kNQc8bo51HKF6XrfJ46Ul6+dnNsvP5njw4AFbu7vkig5JB9oagghh0NvXhdDaibZ10hjyAYL2sEGqXKU52E532GHy/hTb+0kSe5u09w/Vyh6CadLf1wVAOBIkWyjSGA4S29xid3ePpta2OlqT+1sksxlmZmbYTeawC6XqTW883RieGb3C2uwUUw8eki/ZrO8dcLC5wqPHszjSIH6wRWtfPwCtHZ2EAlYdhttbG/SODAPQ3deNALZ2tukf6kdKSXf/MInNrbp+3tjeIrG7yfT0NCXHpFz2DvpBwsDZqyRWHnFvcop0rojApKuztUJPWweNkQDCDGCKAps72/QN9lUU/OAI8c1NdlIpuqqL9Xr6eo70eYWuSn+v7+2xv7HIzMwjHMeoWDNdlajJSKSBzo5KqHbAAkdKenp7MYXA9EfwkSd+sEVb/yBCCKLtvZTi+wD0D/TDMXKIgN6+XixDYAVCSEok9mK0DQzVD1xSspNM0d3ZAkBfvwoKq9xOOg5tDQFA0FOVH7cgSKCxraMin8LA9B3FXP3pGOlvbdzyo8vUO/gsV84NUe9Y9YfUKyxUCOEZbakzoIJJ1HV9iqEzrG9Gqntu9amH8lQX41vsFgN8aOwys3cTOHYZs2yTLZZoCAbIprNYmmc6k0pRluA3BKmCQ8iodpeEc5euIpB889uvMX5xiMTmDnZnA3C485GUFTPdcRz8Ph8ln5/unnYebxzQ393JSFe0TvOGw1E6OyNcHR2sbXy6u/kERx7OY2t96JQplGzCQX8NQ9Mf5ur1MfLpPSanZ4mGwoxeGSMaqES8JreXiO2noaeZXCZDvlCkVCrVMIw2RNlKZ7Fa28hmsti2oCEcZnd7j9aBdhLxDULNrXXRgZFQmKbB03Q2Bise+FKu4mU3DMp2xZzNZ7OUbYlhBbg6doNSPs3NqWlOtZn4/QECgUB1SXQZQ0ik4xANRznYT9Dc1UgmsY8vEiVYzFJ2BIFAgPheHCtUolAoaEcHGkhZCRJqDEc5NXqJxkBlylrO7dcLMCr8WGAaJql0pmKuS5uSbRAOR1nbimN3RvEJG6uhkVAwgCDvKYdCCAxhYIjK1A7HwTQtLH+I+NYOhbYIgUCAks+sbJHg81EoOUQDFomDBGa4Erbv8/sJYCBNC6RDOpGuhI0LB1lVhImDVI0Hn8+HaRhYPj+lUhnbdmrPkx4wpforGAzW6FXnlUgp645frODyzjzLgGNRfY7c6/afZ/Z4aSK3w0uvS93XTRy9vDuf2ynki3bgpO4ycS+FLBh0GHBp9AyTd+7S0BBC+iu+imAojAAiAYOZ+/cROER7hgmYgnAoTDET597ME0zDoKmlnWhbP5GNe0zcu0cw3MipnjABx8QygmBVzDnLH8BnGiTjKQ52d7FzSRZEgI9++EaNj0hbH5GtaSbu7RLwBzl/6TLhcBiBIByOIISgJRBgavoR3VHBpt3CtdPdNf5iy8/Y2EvglEsMDJ2lq2mIqYmb+IMhApFGLpwZxrd2j8n7u4Ckram1DsP2oQus3r7N5N4KwoCWSCvdgwNM3b/HxM4ypRLc+L7xuv46df4Sk5P3WfcHCUWauHhuiEg4jBluxlec597kJE45T6S5h92NZVa29sGxGegfweccQHUaFgo31PoqHInQe+oC9+9NcG/domQLbtwYw3TamJi4y1o4QrZk0G/VhyKLYBsi+YinSyEuXb7E9MQt/IEgwYZmzg22EglVIjV9gRCGWXE4BkORyoheSHF/aopyqcjp0UtEWiJEYlNMTu7i2JLL4zeQzgHh4OECKl0OI+EIEgjXHgpBOBSkoa2PyMZ9Ju9PEoo0MdIdIui3GLpwiYl7E6wGg+QLBv2WoBSMYBmCKxfPM3HrNn6/heOPYgrB8OAg9+7cxW8JHH8IAYTDkcOHMRhCCOhoiDA5Nc3lq9cIWkd39Xq96YP++U49y+Ib3/hG6uzZsw269oLDLc/dr23Un76aTSdMf/+sl9G/Q/16EF3z6c4V5RCVsj48VnO61DntlIPn7r2b3Bj7EEJwpKzbs1wbXbQINr1jLMtC2gX+6s4k33ftWqX+127yysc+hiUOnUCqztfD8Onjh/SdGSVg8J7G0L1a8YUxrF7Xt8APBAK1628GQ8WPU84xMfOED1T75QTDN4/hG32WZ2dnk5ZhGFIxoZtn+kIU/e2G8rLqzCuAdGZVUoQqYvXOUES6N0pVbam6DMOo7UCk4tt1xnR6pJQ0N7dSLBUxxKHTR+8MffqjrusBLQogKdURbxY9jWEeP54FJJ3Dp6luO1BXzxvBcPjMOfz+o8L3XsNQCZ942zCsfFfCrQvlm8VQyaGQPpobG08wfAEM34QcCktKWYvgdO+Qoz51kHWtrCe3meNlJrnvu+vRTSJ1z13WHcOu31dlRs9drHWqnnSBcI8wulCo3zoGp85fqvO/CC2PPkq8LBgq0/XtxFAIUbeYSqfjrWCI4ePc6dMnGL4LcihlZQ9OqYhQhXUA9Ubc8ey62XZc4IgbxOM65o0mL4Cfl9x0KVNML+v+ruPg/gPvLclOMDzB8Hnp/Y6hEAJLSinVrk66KZLPH0bZ6WaPHkPuDgJRDephrfporJt5uimod5Qeu+7WiOpT16zuNfyqfscugVHxOOta1ikXOEjnaWmMks1ma2UbGhpqbem7V+uBMfr6AgWwodX/ljGUDvFkio729qMYOmVyxTLBgO9dx1CPAK3D0HFqvL9VDHO5XG0J9tuC4XtUDt84hg7xZJr+3t7vnhw+B0MppTR080VlVkln7jgNp2syLy3m1uh6veqaWzt7aXl3R0npcHAQ98wDsLc+TyyRO3LPLqZ5urRWo0N3Oum06JGlqrwuPKq82wTU+Uwn4ji8AQyxmV9a8sRQ5reZWVh/hzB8cyOsPvLoGLwVDB/MTCKl5Mnc7HMx1Hl9s3I4/XhGyy95PD0LwMHBwQthmD2IsbqTeFsxNHB4urj4pjB8o3L4IhiqeoQQh6tOvRh0A6dXcpy2dZfX3xm7GfUq7waiWhM729t0dnUhpWRvdweLEt+ZmGH03AVGhvsxjfpj70EiBEi7xML8MkUbhoZH8AN2Mc/TJ7PYwsfw0ABISfJgh9X1LRpbO+nuaKGUS3KQzLO1vc3w6TOIco619Rjhxjb6eztBA1x1QCmfYWUtRqixhf6OJm7dfo3uwTOcGh6pc5ipz3w6weLKOuGGBqjGD2SSB6yubxJtaWegrxs0YTzY2WR7P0FLRzc9Ha3k0wnS+QLb2wecHT2HnUuytBoj0tRKb2fbkT6RUrK/t00mlaaIRW9nK2tr64Qb2+jrbqeQTTG/HsMXijIy1I90bDbWVkllshhWgFNnTpGK75NKJChJk1OnRkBKdjbX2TtI0T98mvaWqOcDt7O5zn48RUfvIJ2tjdVehZaWytZzhWyKhcUVgtEWog0B2pqb2D1IV0LQ7TJ7+3G6u7vY3VxnL56ipaOH9pboc+UwkYzXyWEqmSQd3+WvXrvN6PnLnDk7guEqD5KNlSUO0gWGRkYIGkViu1mS8X2sYAP9PV34gmEaTB+5dJxkJs/B/gHt3b3kk3tkCg4jp04R8B3dqcqxS6wsL5MtlBkcHiEc8JFNHfBsaY1oY5TKzoLeYQdez4zK55bDd+pZNoQQRrlcru3QoxrWzxHQkzpXwTRNQqEQgUCAYLDyHlydu6DMF6UVdU+u+tTNvFwuRy6XqwWbqL9SqVT7W1tZro5iBsvLCzS2tNLa0cbwUB+WtmRX8eL3+7F8PnymSUtHN32dTTx4+ISybbO2tk57dy8tIZh6tADFJHenn9E/OEh6c5759X3yqS1uTT9laHiYoCm5NzlNV28/ud1l5tcqi56Ux7lQKFAsZLl5+x79Q8MUD9ZY3svT1t7M6TNnaIgEj2BoUGZi6hGnzpwlJIpkCxK7kOb+w3mGRk5h5PZ4vLhRUbSOJLG9wtzqHsPDw+wtz7K6m2J/a5GpuXWGR4YopPa4eXeajs4u4hvP2Erkj2BoWRYTEzeJtHbR7Cvx1VcnGRw5xcH6AuliJRitp28AM7/L7PIWm8vzGNEOzp4e4iCeImg4fPvV12hu76Y96mNyehbLMgmEGjh95hSz0/fIlewjRwUaQhAIRhg5NcLczCTZYhnHtkHC0vICUtq8+upNOnp6CcgMr92ZArvEyvJaRdaEzdrGBiCxAmFGTo2w8GQGR5jPlUOol0PHkYQammlpa2R4qB/hIYez9+9wUDAY6O1g4t4kFBN88+Z9Onv6sHLbzMfilLL77CSzJHeXmV3dZ+TUCBOvfh3b30RfVxP3JmdqchgMBvH5fBXz33FobGlnZLCXiXuTlApZbt19wNDIKSw7Szp/eN7HEQyrfBiGQblcrv255fCdepallNLQNdNx04bjNJT7vq7Z3OayV10qKYKeP2VRlgdVITAxDROfCwBVn6hmdqTD1voqy+tbpLJZBNA7OEg0Eqajbxg7s0NsdZGhC1cIBYOcvnyN3aUlQDB85gyhYIBcaov9TImVpUWyJUlyP3FEgxfTu+xnSiwvLpAtOiT2ErXDedx6WkpJPrVDtHuYSDhEz8Aw0bBFYnedzuFzhENBhs5dJLGxXsVAsBHb4NT5c4RCIc5eGGVrZR0QjJw5TTgUJLG3QbYMqyvLFEo2BwepIxgKIWhu76K9OUpHZwe9PV2Eg0Ham8PkikXscoHlpUX2khnSmRyOlNXoRkEwVFF4vYNDNEUjNLd1YNs5QJJJxnn2bIFkJkuxfLiHqkqOdEglDip5sjnKDiBEZbd0AbIYR0S7aGyI0NY9QEdrRWB1iZFV3DLJA+bnq23ZR0fh58khQiCq0yafz1tulmNbFNL7LK2sk0vnsaVkcGSEaCRMz0APqVSyWj8IYTE8MkgwGKKzq5PennaizR2YTvooBo6DlA47mxssLK2SyRfIpysy0BAO0dNfkQGdH3d5fYMb3RLX871Tz7IQonIwstv0eZ45o5s7ugPJa46jN6QT70WkVwcfXneQKA9tiXyu+i76GLCklEhACIOJiQmujH8Qv2GzOzGDBPL5ylbsODaOtIiEIxxkstDUhF3IIAOVB8MyK5rctAJ0dfdy4cLpug6pM91MH51d3Vy8eLF2/c7tlSovR19FGaaPcqES/uvYZUolm0AwTCGeBZqxS3mkdXjqVcjvp1AoIRqDlAs5jEAAIQqY1UhKvy9IZ3cDZ4e7Kvssan2j95eKPVFUKT6ccoHpJwvcGB8jn1hnbg/6Bvq5PTVLvruLa1cvgSxiqtd61Qdme+kJGaOVCxeGyWcTdbyqNndX5sgYLYyODpNNV/wFqm0kYPiQpepxi9KhkKvEAjiyerhvuUipaLO9NEvaaK3WU1nzoaa5XnIoSg4OYAqBXcwifYHawOMlZwDhSCOnTp8hEgpy4YKA/CaGqL5mdGR1+nnYnjoKQEh5CCr1z4mSkenJCYYujtMUDhDb+SsM04ddyNRkoFzSNmVxYai/TtUtDrccvlPPspQSy7ZtRwV/6N5X/cwOPbDEa02HEIdRZWo6IISoTUHU9+McYeFwuNaW7lVWbRqGRcAS3Lk7gbRLlE0Lw/QjcmkePpnn0oVzmELU+QWUGdXS1MCDqfv4LAMwkBIKyQOmpqYoFwsMnbtIR0cDizdfYyIWJpvJcvH6DQqZNYr5fOVot1ALgfIC9x9kMIXB6fMXiYYOwfX5fPibe2g01rl1+w6mYXD6/AW6WlqYun+fi5cuE/YZdRgGo51Y+QUm72fBKREMRwm39FBenODuRIxiPs/5qzew7ThISc/QGe7cvctOQ5Rcrsj4K68QX3uIlBWMOwfOsnbnFk/mEkhHcu7iJcJ+S8NQ7eJd9Z6LynkZyuQ0LB8WRR7PPkaW84SbByhkM2RyeVLxfabiKa5eHEHWXqtVHpSG5hZmZ56RP9gknswjHQcp64OXgg2NbD6aJ7O7TipTwjQMTMtCVh90YUXpCNs8mJ6p7LjumNiYyHySqQcPsAtZhL+BYEOU2ONKPcl0EQHcuXmLD/3ARzGrD44uh2dH+vjOt79DOBwik0px9tK1ynF+jsPkgxkuXrqI6ZLDaxfPMj0zQ9DvI9LUxukuC8OorrswK0cDO46k4hMztHtW9aGWtaMClRwqehoawjyemSbgM5H48EfaMXOLTN7PIO0i/mCkbuNcHUP9DYi+5Fx3aCr5fyeeZUCIb3zjG4nR0dFGJVA6cfr2XgpQ1bAiWmmeXC5Xe2WkKwX12gbqQ1PdR92r9vU9GhQ4uoJRczC3xlR0q0/VlmFUDl9R9amtyBSPNeeTBro72k/vJC8HlP77ZcLw9t2bfP9HPoZpGEx851v0jF6nJex7xzG8PXGLD7/ykZcCw5dFDh89epS0DKOyWZY+0rtT/VuGo28uFHHuOtz51Xe9nHtepZs9enkvcNymlbs9L1+JHsjiRd/zktvc0zv4ZcSwIxrl3r17lZPfzDCNIatGp8rzTmDo9/nrHhqV3o8YerWl6FT33g9yaNs2lpTS0LWNKqh7id0HnyhNqXeorq3T6XTFNHPl0V+h6nHv+ntk/bq+XF335OqmmttrrMqqzVeFEHXBJ7pW1jtRj8/3WvCj6lE8uBfw6J30smA4cv5S7Voul8MulbDfBQwvXbhMsVh8KTB8WeRQCCEMx3Gkrp0UQbr2cSd3mKlq3F1e/+0243SGdOeK6jS9Hn1RzBtJXvQpJ5GeVP36SOJOXhpXXXePNCcYnmD4evS9XzEUQgjDHe7qNm/01256ZV6AqevHhdC6zUKv+rzqdXeizoj7uk6DO5+7bp0etyAdB64XDm6z7nsJw0I+j5TfSxhKyraNdGxsu35/Fr3cSyiH0pJS2upIs0KhUNNa7nMH3I4eIURdPLmu4fTzFHTidDPP6ywDNzBeb0+g3lQzDIOFxQVGhkeOtItTYmE1xvBAf11b7vp0XvSOUFioEUXflahQONzOXu0dsLC4QF9ff+314tuJ4eLSIqdGTr1jGJbyWfCHCHj0nZSVNwVeGD6YvsvotQ8RNN8eDJ8nh4vP5ugdOk0xm8VqbPTEMJ/N4AtFMJCsrK5w+lT96254MTm0C3EezG9xdaiRmY0yY+cHaxiq5CX/z8Pw7ZbDd+JZFkLIyvHNHDVn9MrclSjA3Q3qeb0CSPT6vTSfF3jqWjabYW9ni/14inKxwMb6OulcZT7YGI0CkMmk2d/ZYj22hSMBYRBtiODYJTKZDLH1NZLpLMV8ho2NDUp2/eijUj6bpfJKXWKXCuSLZQQOmxvrJNOV10q5bIZcJsX6+gb5YgXoaLQBQwjKxQKxjXUOEuk3gKFkf3ebrZ19crksssqHwjCdTlX2bazyWMilWVtbI5nJeWPolEhnsmzFNtg7SEL1fiGXYX19nWy+skGKY9vsbMXYiG1RKpWYmrjNs+U1svkSmUyag71t9g4SZFKpWjxLNp2iXO3XCs17CHF0tFJJCEEqsU9saweJIJ9JU90OlVRKxZiUiG1skMrma32YTsbZ3q3EY+QyKdbW1sjkCkQaojjFPK/dusnK6jol26n2wTrpbB5pl7h75xZLq2sUSjbRaEMlmMkusRmr9AeAwCGTybK9GWNnL368HDo2mUwlqhjpkM5kEEDZtgGHcjUALRnfY30jRqlqaWQyaXa3N9ndT2CXi6yvrZHJF2v9v7u9yUZsq4KlY7O1GSOezByLof48uKcw6rqiWefj7XyWAWHIag73A+0lADoB+onoXmaMW5Mr5eEmxKsNLwa/8dU/I1N02FyY4cvfuoUwLe7cvEXJkSwuPwPgq1/5Y/YzRWQhyZ3Jmcq6kOVlZDHFn33lqziGxaN7r3Lz/hMsy+DWrTvYHpFxhdQ2T1cqZ3MsP31MulDk9q1b2MJk/uEEG/sZpu99h9mlDfw+g5uv3cSRsLj0DAkc7O0gLD9Ls/fZSRWO8Kdj+HTmHrH9NE4hxZ9/+SsUHcnszEw1Lzx+NA3AwtI8dv6A79yZJhDwk4jHPYPSnNwOf/YX38QWJluLD1naTJBP7XLr3gw+n8XDe7fZSxd4PH2HRN4Bu0AmV0SYkoZoA5ZpcPNbXyG2l8ayLJ7OTNXOYnk2O01RwvzDSTYPMjjFDPOLG56Dg2EYxBZnebq6DeUst+89QDgFJiZnyCZ2eLKwhlMucPPmbYRp8XDyFvuZIhM3v87y5j5+n8V+bJEHc8v4/X6KxSKrK8+whYEwK4rZNAT7u3v4/X7u37lF3gbDgmhDFNMwWFyaB6fMa69+B0dYbC3P8fjZGk4xyZ99+SsUHUFia5HZpU1POXTKeeaeLlQeLrvA7JM5cMm6Uy6yu5fAb0pu350E4Gt/+SXSBZvYs2n+/Ju3EKbJ7dduUnIcpu/d4iBTxMChXC5x89XvYGOytfyER/OrRzB0TxO8njmvQVmXtbfjWQakJUQ1KMeoLJX1cr7oZpi+/FaZN4ZhkM/n6xwvcLjJhyJCP/1ZXyrrDibRQVDXm7t6GR7oo9Rok14p0tbaQltIUJCHdDZ39TEy0AvA6vatmgA7UtI7NEJXRztOop1Sy2m62qOsLy5QLNtYov79drS9j8cTUzgDbSTzkgErSyIviO/vYfl8LC+u4Qs3cPHCeYKmYHdnA1scxu03NDayvrEJOOwlc3Q1hY7FcCdd4qMfOYtpGqytLVO/I3g1wMyoBE9ZgQaCosR+IsvQQO9hNKWGoeOzGDp7nt7uLrqbBPcWdyjJfUavjtPRYNES8TH9bI3upmZWYhucOn2alqYGwuEwjU3NmAZYja2cOz2EIQSOrJrtUi39d9hO5fnI5REE0LeyiF0uY5viyBuHx/OLdPcPUyhJkvsHRNs/QPvuDl+9Oc3Hf/hjJDefkrV9pJIJgn6T9Vgcs6GFc6eHsAyDW49ifP9Hf7B2jsaSMLD8ASINYVpbWxFImpqbiG3vIJ0SRSNIMBiksakRU1Rwyae2CbQNM9DXC71dvPrqBKWeED1Dp+jqaMPfGeHWo1Wg54gcVr675vSCyqbBVHadLzuSgN8gkcqSrgZRNXf0MNDbTSlSJLPu0NnRwd7yPJl8hmQ5wKWBXoQQ5BIbBDuG6Wxvpau9mZs373F6oLMOQ/VQBwKB2vRJ7ablfg2q5OqdeJaFEKK2Ya+edG3mNll0RnTzReXX50NCHN2kV93zak/XhPpqVQCfFglnCuWsqVf0fn1+rrVjCIGlgAfM6qavCKph4fVzQ2GYtIUM1lYXCbYNIIC2wCmuugAAIABJREFUzh6GhwcAsCwfD+5vHa5YNIwaiE4xw517j7h67QrFgEP8dTAUgiofshYdqehCOpSL5VrYM4afVz78EZL7O3z7tdv82A9/rBZcrdqQUtYW1qnrhqGfnG2DYdDVP0RHT5lnT6bZSfTWgBRC4LcsPWgbWXVglotlqGIoNPA9MRQCfyjC0NAQAb+foaFhBJJsrkDYJ8iXKiZ8V28/gwNthMOjGKbJ3YnFw7YdWV2foo2e1f8CyOyvMbN4wNULZyikdo/KYXUqStV6RDrIquLxqdFUiFqtR+SQQ3msLO5yDikQAilhafYBTrSHwYFBNnZ2jsqqoSiWCEPgOPouVyY4hdpv6YFhrRdcUwx38pp66Dy5+XPL4es9ywCWlFLoFeuvh44zYfQKDhn33pHYzcDhdvtHX8/ojLjr09tEo0enTM8t9GxCewWEwNHpkip8t/6BGxwZ4o/+w7f5z37up/FRRqbnWFkzsAR09PRXLRbncCqgLXSz7SJ7O1vsra/RdKabJ5O36RgdpyVooicpJT3NER48miMaEKxvJ7gqIRSwePJ0AcPOsXmQrtQtBMV0gvnVGH5LrfE4iqFdowRENRS5f/gMt+9PkOvtZnN9nYvjHyS2ukTBFpRtiYmgIdLAwvwzzo4M1tXZ3tHMzMwsTSHB4voWo0LQ2xxh+uEs0ZDF1m6ay3BE2KSUnO7vYvrRHP3d7TjCotEs4IS7+IELbdyenOLG9QukF+6yZhYJWCa9QyOVOhyJg8PZoR5euzVBf1crkcbmamcLQkIwv7RMa1hQyOfYiq0R29yja1QSDQRZWFhkqL8fBIQaO7FTr/FsQZJN7NDZP3TYd1LWy4xLDoUvQDGXZHFpieRujLztr5M3ISoDUSqdYq2QJJUuHJHDmoQKgTBDtPhLPHzylJBl0NM/gJOaZ36hTD6xT0fvwBEM9d+65aZP8d0+C/X9bX+WVbi324PqDi+taT+tYuXRVZaA2xxSzKi69CmGHiqrx67rppMe7loulwkGg+CUSWWLBAM+Cvkclj9IqZgnEAhW4v6rb3ay2SyBgJ9CoUgoGKBQsvH7LOxSEWlY+CyTQj6PLxBAUL+bs+Ijl8vj9/uqtJQpFUtgmDQ1NpLJpPAHggjALpex/H5KxQISgVMqkskViEYjIEweTE3yygc/VLNE3BhmUklsYbL4dIbRq68QMCSZTAZh+vH7DCzLV1nuHPATj8cp25KGaJRgwH8UQ6dMyREE/D6QNtl8+f9v79ua4ziSc7/q7rkDA4AAwTupC3clQiQlL28ipXX4PJw4cfxP/Hv84H/hp3PW4TixjpXXsiRKoiiKK1KkeAdAggCBuV+7u/zQk4NvktWg1rvaI812RUzMTHdVVuZX1dlZWVlVKOQDhMM+Ot0+KjNVFPIB2q0G2p0e/Fwes5UyYC0ajTpKM1UgDlEslsb4t5p1WBOgVMgjyCcPTKvZQAwf5VIevp+DMW4M+90OWt0eSqXE0Tw3Pw8DoN/rw/gejI3RaDQR5IuYmSmPMZQhlvBdKleQCzwUCiXYOMROrY7ZuTmEvS46/RAz5SK8XB4mDtFoNFCaqcLDaB2FjbFTqyFXKGOmXEQ4HKA/jFDI5xD4HnqDIfK0noP7YRQOsVOro1SuJMdMlIvoDUIU8x6a7T6KhRwatRpMroB84COfz4/7IWyE7iBCIRdg0O8hXyzDMxbNRh1hbFCtzsIzQKNeh58volIqOjHkZyGO4/FaKh6S8HP3YzzLt2/fbprf/e539ZWVlaq1dmIahmPLOW6cLQXeVmzS7H15OzOdn3ci5sU2TJ/fVrxIjHdA5rTXVuuSdLSa3GPQ2UEkY9c4jhNlNUp8nRfkvIwh0Ol0Ua1WX4nhN9ev4q2zl5D3MgyzfvjTwvDWrVuNAICRt78OIOGCaeMh/duYybMPeBYkbbzloue6x2bZXvddvHI+l2Z1ycr3GUD+L5jthaGc6vQqDE+/ex7G2AzDrB9O/P+pYBgYY0xyBF00MXPhOjRFQJc8HNjDArBgPJTg1XUsDAeEcL3MjyzXlTzMgySOjefOwIDLWQ/GTB4Dx28DvSEq88L0+W0gsv5pGPoZhlk//EliaG1yFMD4gmTizC4tqQntdc1VqV5RmKah5dsVOMVl9IwL52VQdT26Qwm/HDOg63xVXZr3DMOXecow/PlhCACevsEFeB6X72mBuWLWnsbsRpyxJtPCaMakHAt589sbTmCvX/sUQ7zaXAN23yIvnq+jH04GiaU1itx/+uxp4tHmBo1DPN14/tIaBI2hjCv3wvCbm9dhR/X8UAxt2MfTzRc/GEMX3roT/1AMAUyY9j8EQ34T6g77Kgy53JdffT6erv1L98P/LoZDdTLZ/28M/9hnGQACY0wsZgrvliMmjTFmvFGH1kY6xl6cNuKAsdZOmFv9fn9Mg01BNr1YCDHnkgdumJhTcZxsPpvLJUFDUYRwMEAYRShXyuNt45LQaQ/5XLJRaTRa/NNqdxBFowcYNglA8QPkc7udKckbYzAcolKZgecZFAp5BL6fzIoMB4hiIOcDxkwuZzbGjDc67Xa7MDbE13+4g7dOvpnsYzmSPwpDDMMQhWIRge+j0+2MTcQwDFEoFBKPth+MNlX1EMd2vHlJFEUo5pM9SM0oFiKKhvD84CUMAYtut4dyZQYeLKJ4dHZGHCGMkWwJN+I/8H0MwwjFYh5RFCGOIvQHA5RK5XF8ipypGUch+v0h8oU8fM/DcNBHZIHCaCen4XCIKAoRBHnkcgEGI3kSWWIMhwPEMZDP5xDHETw/mZ0IggDhcIAonnQUdzsdGD9AFCVxE2b0EA5HeBnVD33PQzRy6iUzY314flLXeLPeOEIMD4V8Dr7vIRyGCKMo4dMzgI3RbLVRKBQBWBQLhWRzmFx+zFsYRjAmmYYPo2h0unyI4TCE5/vwPYNrf/gGZ8+8Oz4IWTDUD65+DkSZ6PUm0td4+blrWPTnepZ938fLu5Zib3NMP9BpWtFlAon20+afDsDSie89vn8XvQjY2NjClb/9EMNeEze++QNmiwG2m118eOV9PPrua2y1Y+QRIQwqOP/uKfz+3/4PZhZPYHFpP+obD/DawgF8+8WnKFcXEUUWb6+cQn7Uia998ltExf2olnKotQb48MoFPHj4PfYvzuPjjz/D0v5lhLHBW28cwcMnT3D44MERfxZfXr2Ki5evwFqLr659jrfffA3rz9YxPzeP40cPI4HK4tG9uxjCYHunicuXL41AAx4+uoelxUV8/cXHQGEOCHtY3W7jf//6PK7/4R7eWXkLJu7j+jff4f13T+LBk6dYLHTwz/96Dad/+TpatS0c+uV7OLE8N6IZ4csvPkd5dh71nR28e/4Cbl77Eucuf4D7N69h6bV3sG9mNN1c28A3369hfqaI9sDg3LuncP/ubUTwsbldx4cfXB7v+VnfXMWdJy8wWy5g6cARtDYfYacH5E2EoVfG35z+JT767f/F4uE3YXtN7HRiHD64hBdb27h45Qqu/vtvUJ4/ChN2sLHdwfFjh7CztYUzF66gt/U9Hm91UMl7aHRjXDr/Lr6/+RVedC2KPrD2vIbzMLj77VfoxnkEdgCvvIjTb70+7nOP791CY+ChlPNx7I1f4MG3XyLOzyLutZCrHsRbJxbxL7/5DX7x1mmEvSbKiydwoDLAje83sFgtY2ZhP44uVfDpF1+jWp3Fdq2N99+/gK8+/ximOAcT9rFW6+B/fXgON775Hu+9dxqIerh+4zbev3geD+58hxAenm1u4+KvzuDZs3XsW1jGiddPoBDs+qZYWXB/lyUSLuuOk76vn6E/57McaLNKZ9JMusY/f0xyMZFmgrmuHzn+GpqtNtq152j0Ytggj9Nnz6IcGDy4eQ2b9SbWtnu4cuk8AODTj/8Tw9gizs/g3K/eQzgcorlxH0DSKJXZeRw5dACBR+HK+SLOnD2LUmBw88bn6Ed2ZBAkQV37lg5gvlqBsYNR2C+F3dpJfmfn92H/8jJOjMLQE3mAY6+/jnqjhXptB73RLtUSv2PDNhphBb8+fxpAjJ2PPkpuWsLN7gYUWWtx6MSbWFl5C3E0wGeffYUTy5cBAI3NJ+ibWRxfXETFH+LBag1/c/Zt/P7f/h8OnHgb++fK47fT19/cwhsrZ1HwPVy7dgNhfAon3ngTzVYbO7Vt9CKLipeY5ncerOHC+5eBOAZsiDt3uvjg/Yuw1uLqJ58igkFudh5n31mBGTbw6bdrWDl1Cmt3bqDW7sMUZ3Hm9Aq8qI///OomVk6dQm3tDja3G9hc3cSVDz6EAfD11U/Q6PTwrD7ApQu/AmCxXduGjXvYagOXL6wgCAJ88vEniEfKAjbC2mYL/+Pvfp1gFbZQH5bx63OnAQAf/e7fYY8vYm75CM6cfgc27OGzr7/FodllGOPh0LET2Dc3i3s3P0f1wHEsln10a1vYeLGFVjSDD06/A9gYO//x+6Qxx/00aaI4tjj+xhtotTrY2nqOMChjaf8STp58A6OAzolQbp1cUc+u50Xy8tSoHn5w2T/1WQ48L2E/bbGXCCaJ52NzudyYQdaCYmIJA1oYa+1EfDszzfsCsuc3jmN0G8/x5c2HePP148meAgB8z08ObLUWQIx+v49o5Cew1gKRHZmpeYTDIYrFIoJcgHw+j3MXr2Dz2TqufvoJzpy/hNlCYmgFfgB/dEx6FMUYDIaIogiR9XHp0gWsrz7GJ7e+xcVzZ8EhfXEcIxoNkwwsojBCbEchy4Rh7fljfPdkB0cOLI3uJZsLe6MVnD4ixJ4/xsgPkjBhGXvaMEIUJqseoyjCYDgEkGAaxzE8Q9GUcYhgFKhWqC5jeWEeHgaI+l3k8rumrbUWEYBhv4fYGJxaeRuN549x+/ELHD20jMGgj+EwxBAmMU2DAMVCAcPBALAxfJ49QGL+y3L34XAI3yTfNk7OxAh8PwmnhkV+bDIDNo4RWotwZDr7xkM4HCL2dv0OuUIONo5g/KRcLpdDYJJNgDEK60Yu2O2Hwy6sRyd7xckQpJALEp6iCGEUIj+zhPdWKnj44Ds8CGZRCZPNhY0xOHZyBYvVAA9G+1laa5HL++rBjRBHMbafPsCtxzs4dmg/+oN+MhyLY0RRiHiENQ/VhU/P8yZ20+KHXQdf8fOlFc6P8Sxba5OSfNM1bmJnBzPG5Vg41m68ck6bXDIs0XPC7LzZrc9g2GvD5MsoFQLUduqABaJeF3fvP0KzvoNHLzrYP1dFNRji4dpG4sj0A+S93RDoXQ9zjKdrT1GaqaLsx+gOJuuCJRMNiU0RDXp4tvEC1YVF2EEPUWzHlkSChYfBoItao4lH925jux3B8wIM2m202h3EI3l6rSbylSqKeQ+1eiORlRrUFBZgmhvYrjWw/ugutpsRTJBHs7mDRrOFB/e+Q7u/G67sGYPVB/dRazTx4PYNzB85OcZwfvkYho3nKJQqyPkGxjO4fv0GPviff4/uxn3U2rtj55NHD+LZVgOVmQpggH474bOUM6g3WhPtfmxfBddvfY9mo45WN8ScH+LR+nNsPltFzwuQJ4eiMWZXqRoDQL9NqW8Z4MBsAXcfrWPnxQaet/qYm62gFPWwtrGFrWereLbZAvwSSnETaxsvsP7oe9hSBeNHyASoegPcX32WWG62glx/C083t/Hk/m3kqgvwPDNRvzEG3WYdjU4fS/uX0W40cPy1N7G18RSlchkGFn5pEabxDC9G7bJVHwJ+Dq3GDmqNBu7duYV236LfaaEwU0UhZ9BotGAM4IURdupNhKNl7PJA6+dFP0f8zc9I2vDix3qWjTEwH330UWNlZWVWF9ZMCIPsb9D7/2mBgN3xFzssxdrQZpBoXO2RNcbgxYstLCwsYOvZOjqhhwOLc/CLFfQ7TYSDLja3mzhy9BiK+UTzb6w/QT/2cfjwQRRyOdRqO5ibm0ehUECjto2Z+UVsrD7ETqONxeVDmJvZDZxqNmqozM7BMwa12jYqs3NoNupYXFjAs/U1tHtD7D94GLOlHHYaTSyOjuCz1mLQ6+DJ6hpmF/YjH1jMVefRqm9js9bGieNHx6sVnz9dQy9OjhDMlypot+oolyqoN2qYq84jCvtYXV1HubqIRw9v48K5Sxj22njwaBULS8sIfIO52TLqrT6qfgNf3m9jecZHcXYBxw4fmMBw2O9idXUNCIo4cnAJjXYP+xcXEIV9NFoDzI5kBywaOy/w/EUN84vLWKhWsLWR4H1wcR75cgW+wXgFZH17E083d3DoyFHMlPJYf/II/djH0SOH4XsGtfoO5ucWEA37aHT6mJudQdjvwOQr6LYbmJ2twiDGTr2JxX37EPbbGCCPUs7H5sY6mr0Ix44dRc73ABtj7cljxEEJ89UKyqUSbBzh6doq/OIsjhw+AN/zqB9abKyvojOIcfTYceR9YPXJY3jFWSwtJKHgjVYbC/PzsHGEequNmWIeq2triBHgzZMnEXhAr93Ak7VnKFcXcOjAEgbdNtbW1lGq7sPjx3fx/oXL6HeaePhkHfuWluF7wOxMBZtP19GJPCzOzaBYmYEddrH29DkOHT2OYs6f2PWb9+nksGtO/Nxx/AVbAxzB+ed+liXcu3bmzJk5ABOMynSfDAe011RCRyWxx9W1zDzNV2Ht7s4/woMWWOiKcGyGSb0ClqbP/63dnZ3hstrhwxp/7PmP43Ekps7PIcM/BoZXv/wMF89dSsUwaq/j5lPg4juvZxj+BfvhF9eu4tKFy38VGN69e7flaRNor8RCaxNHmzmS9CyHaFOXycN1uHYE4mtpGlIPdzRtXS/LojsHNzYPp9I63A9J/x0MT586syeGpriEd944PEFL4yXprxXDH6Mfnn7n7F8Xhjx20swxUU2QGdbMazCkUVzgaWZd5lOaWcUNovlMM8O4QXUQi0tODubh65rnHxPDSqWyJ4YwAWbKu4uLMgz/Mv2wUq5MlJ12DANjjOGVa5KJTRr+zaYdn5ugV9DJh5ers+nLMerMtNAyJgkm8X0/CUCi4BCOiExL2tySOph/XrorDcZxIHEco1KpjO+32+1xWd5ViZcVZxhmGE4jhgCsZ0eb3+xlxqRpar7HZfcyk9hsYwC5PDeya85Z85CmHdPk0fmlcZgv15tHy6PfGhmGGYbTiqExybZ6E4zrgi5mXEkDrM0gfY0B2mu6hxuV4zT01mNp2p3rkaSDVzRQXL+rI2l6+p6mmWGYYfhzx9Bai8AYY/V4SIJDJLGJIt9xHE8ETbHQvu9PeFpd2pzrZG+w69BaYNJk4sAVXn7LgPAmH+IZlrh4qZdPeBdvsLW7wWDW2vExehIPMl53oALGND4ZhhmG04QhgNhjzaG1nCSX9jPGfYaBaF75LeW12cf50xw82pTT/OjG0UEu+u2ir3GD6TeMfutwPubTVT7DMMNw2jA0xphAA8AZ2TnD+VgjcWNoplxlGFT9XwDiMjzlpcHSJqBLSBcvLpn0W0eSnnLTncLVIEwzwzDDMI2XnxOGADCxrZ6OFRfi+qg7SWy2MWBsZgltF5OiBfkMEf5mTy8fLcemGr8NOBCFo+L03LSW0fM8NBqNiWW5wgdHxXGwDe+YFIzWC2QYZhhOK4bWJjtlWdZarD3ls5fWketcjivTGpEbSL55PKlNJM0XX3fdk/9sbmmZpPNonuTjKq9NPC4HvHyydYZhhuE0YQgA47NO2bTSIOrxDIPEAmlTSAsk9Jm2BoMbjPPLNR3M4hJSl0/jme9rfl2dgseQaZ0gwzDDcBoxNMYgwMiyEABcTPNn91i3lxvDBa54bkWruQTiXYM4QIV5cplVmmf29LJ3l01BHbcvILGpyeM7jqtnQF0ma4ZhhuG0YgjAeFwJF9RaSTOjiWsPMDeUZoiTnmt2aVptqrmSCwyWRWv/tDeK1uRMQ/PFuGUYZhgyH9OGITA6GFln5v8cdqoZcjHvMsM0KK58rDVdZV3gcHJ1BF2nnqLSMmsaDDLX7eIzwzDDcJoxBGACAIbNGtYurGUksXnDm4hqE0gSm08MNm80KoEf2gSSvHEcT2z8S7v3TAS9iPfYmMlNSiWPbgjmOU3juxpD8yAb9GYYZhhOK4bWWutpxl1azfVfaZ2JpO8ZsxvzrrWkqwE1WEyTG5Pp78WPBiCN9l6ya62s6WUYZhhOM4bWJuHer8zsAlYzq7UZM6Q1pDSarkcLn0ZHHD8MnH4b7EVLrmuPNssp89VcxsUzl8kwzDCcVgyNMbtHAXDAiGTQIEjsuuSR4BPP8yaOftOeXmZGyjIdMdXEYy35NHDCAweWtNvtcT7mYWJ+mDzbvDyZj7STABvhRxpRgmGYvjbphL8MwwzDacUQoBPJWNPINR7TaI2kGeT/+h6bO666uHFctDUorD05co6BYZ7HwqrpsDSZ9FtJwNV5mJcMwwzDacYQSMK9JyqUxFqIAWSCujKXoNxALgFddKSMyyHDGpKnuzRYaTy7QNDlmbbwx7TS5NWyZBhmGE4LhtZaG0ghY3Z33wYmNyxlL65rI1D2ErOgQteYl0NvXYExLIyYQ7qRrbUTxxpyUIrwxh2EtarQdTWSnDOiG4xpsonINDnwJsMww3BaMRw7OF1gMNBa86RpojTtyXWklddx7WlvA60ZhUde5KNlSNOgkt9lprEMWjvrlGGYYTjNGBqjlqhrLegav3Fe+XblcwGpG0ozpYHie0yfQdL3XR0hbe6a87toah4lb9q4kfNlGGYYah5+zhham0ydGmvt+ORuNns048BkrDsHcnDghwSHAJjwpjIYPM4Tk0mYEh54c1G+5zrfQQSVOmRnIfH6Sur1ehNlmC+hyTzrQ190XdygGYYZhtOKoed5mLBjXKaVS7PpvFye82jhOB/TZ23P4O2lVTmvvsa8ac+z5iWNRy2PNkEl8ZhX45JhmGE4TRh6dnRVM5iW4jiemBfWWlhXyBpZfzM4WvPtxU9ana76GERrJ+fMuVG5buaPO5C8Ibg+LpNhuFs385dh+PPHEEjODXkpo97Uk8dwEigiDAvzYtKIh1kE1EEjkvSmpWOGyPTishzEwk4ezs/nJrBc4xPVMRkDz8Et3EnSTD7erJXPgxQzNcMww3BaMQQSy8K4NKg2SzixFuRv1oKcl3+7NOkP0Yi6PheILrNqL9ouGV35XWYa5+FO+Sr6XDbDMMMwTcafIoaBtdayhnQJrSvUAPA1cYpo4YwxToeONrO0YKzdXEKL9tTBJmNtqKaXXHlcMooHWQOa1ugZhi/LmGE4XRiOZ0M0ABKLDmDCS8xajL27/X5/fE9MsjQQZPzGNJmurgdIzDaOmLN297h6ycuCsbnIMfwcA88N4Oo4DJbOq98guhEyDDMMpwlDALuzIVyxNkfYLNH59X8Gn8ul0dH3hZauQ99Li7t3aUpdVxrArjJp9WmsMgwzDKcZQyAZhqQyJlpTH+6qta0GQWvstHwuRtkho8vwt77u4p+F1qG2eqqJaXF5bdaJ3Lw82dXAGYYZhtOEobUW47Uh1lrnGI+vG7O7bFZHenGj8O5D8h3H8cT5Ba4gEYnDlySC6YZmrccBJGxKMdCdTmdcJp/PvxTRJjxzI0pZvS5A6iqXy+P/TD/DMMNwGjG01hqPhWFQ064x6C7N+0PKpplBLBg3iisG3mU6aecS18V5pR4211xmF+cVmvpNpd9OGYYZhtOKYcBMcOLrewWqaBC0kLx6T9/jhtGanvPyfRcIDJrkkUZmYPnN4QJMvtkhpPHQMvDbK8Mww3BaMTRGnRvCQSCuJbHW2rE32PO8iYAWjsN3MauZY9A5KEWDLomnrpg38dZKJ9B1Cs/GTC6oETpS32AwgO/7iKJofAycpsubvvJGqSxXhmGG4ZRiaMenqGvhJLm0D2tpyeMqqxvI9c31MLC6bpcZ5yrzKpp/Cl/6N/OYYZhhmFb3tGA44eBkE0004F4A6E0+XM4f1qBsDnE+138Gl/O46nA1hL4uQGlNzWanfLvkZXOS69ce9wzDDMNpxBBIfBYT54bITdemoNba8dkKkoe1FX8zTRGchXEFinBZrY11WbnOwS163CY0XU4qkUHycLBN2rSZeJJ5TOr7/kSMfYZhhuE0YmiMMV5SbtKkEWL8rQXXeV1lXbS0YtJJg8wCcB4NCJfVZfRv+eg3AJdLk0nn07QyDDMMpxFDay0Cz/OM1qBplWnN5PIYu5hyCccalR0+/M1zzhpoNu9exTPwsiYXb7N+W3AjuqaUdN2642UYZhhOI4bGGARxHBtrJ88RACY9okyA179zgAebOnzuAB+pxtFjevmtjLm4Xq6L4+q1dhWQmB+5J1Fucr3b7Y6vyzJhz/MmOgefH8FypSXpTBmGGYbTiiEAE6RVrjVMWh7X77Q8fI3Hb1rbyzWtaV100lYQMl3Ni9b2/H+vt4SmKW+itJRh6OY/w/BniWG6stirMi4jJhIDKoy7NC//F1qu4BStCbWwQiMNJFfDpl0Ty8oln24UDWpaB9IpwzDD8FXXfuIY2iCOY8teYl1QGJXEYxs2eySPmEAMADMoYPCSW57m4YATpsN5xDwTE07T5jcEgw9MLtcV77ELcKHJZzSI6WitRaFQmJArwzDDcJoxNMbEY8viVebYXoKkmVtShsvqtJd5pn/ztTQeua4004uBdc2X/5DEWGQYZhj+NWAYMMMuYZioMCFjJGGC74kpxdfTzC7X77RGYxNNN7wWmsHX9Qhf/FsHwLgank0y5olThmGG4bRiCACB53njtSE6YEMYZjOJd85hr7JWOmzKCAPazBMw2RT0fX8i2k6u9Xq9MR2JsWewBEQpNxwOJ3hxNYrv+2NPsZiULDsweRQdnx+hA2IkZRhmGE4rhh4Ao4WQ5DKj9DUBXu5xPklao2utyonfAkzHpUHlvvDAGp87hOZDvwFcMrrkSTMVmUaGYYbhNGJorU027NWAspOEzR4xSySFYTixyQY3AFeqwdIgpwnO3zq57ruO80qAAAACCklEQVTK83XhhTsBMBmYIzKKRuYGdTWAgKw7Q4ZhhuE0YWjMaIm6xIizd7TX640J6TMOhLkoisZx8OwNZuFcQgnTAgqPsdjc0uNM+eYpHv4tZpXruDbtJRYZhWa5XAaQmGYSiBLH8QSgvBZAvxnElM0wzDCcRgyttdYTZiRps4SvS+UafAbDZUbxfzbNuEya5tZltdnGvOnfuryWlSPmmA/5r6e7GAPdUBmGGYbTjmFgjDF6zlmbb67vV10TpkTLaW0q90VABknqd3mSmTaDZMzuXLF+m2hwgZfnwtk77JLP1SEksebPMMwwnFYMA2utJ5UUCoWXKtOJNZT2vmqAXFpRKmZTic8y4OATNv/0uQkuDc88yCnSDKxueDZBOU6egeOPjqUXuhyck2GYYTiNGFprrRdF0ZAZc3lvdWKNk3Zfmz9/jKkm94TZtPpdpqbrrcEfzq+1aVqd2pzjt4+rzgzDDMNpwzCO40Fw7969fwzD8B+MMfmZmRkzImx6vV7secny3EKhMFZBURTFxiSnmEVRFAuThULBl9+e51mpKIoizxhjR/csMA4EMcJIq9WKPM8zcRyjUqmMT3a3o3NYoyiyuVzOEDhj+iMnjQUmHDbG9307SmPeRvwzuFZoBkFgSBaTkDd2MBhIdej3+7GAm8vlzOiNY8MwlLI2wzDDcNowjKJoePv27X/6LwuwkpRpxtwQAAAAAElFTkSuQmCC"}]}