{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(to bottom, #3689e6 0%, #4d158a 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/black-linen.png" , "items": [ {"x": 385,"y": 750,"w": 715,"h": 220,"type":"text","text": "Subtitle ","font": "open sans","color": "#64baff","font-size": 21, "font-style":"light italic", "justification": 1 }, {"x": 89,"y": 439,"w": 1322,"h": 403,"type":"text","text": "Amazing Hipster","font": "open sans","color": "#f4f4f4","font-size": 28, "font-style":"regular", "justification": 1 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nGy9e9hvWVEe+Nba+/tON93NpRuQi8BgAEUEoY3gJYKigIhBdMwYn0RxJHEyqPEy6mNGIsmTGMd5BKMZMYiOEjM4qMAocr+qQW7NRbmEICrN/dZN38853/fbq+aPet+q2l/ng9PnO7/L3mvVqlX11lu1atuDnvyzb8Kld74a7gDcYMPhjrmdwgBgDAAGwGFjAQC4TxgGAIfPDbABM4PPA2ys8O0Qn1mOAJ98f8B9A2AwM4cZ5ulFs+XIfTu1uPCELccOg8EdMIPPDQYDxgL4Bthw3w7xeQC2HsO3A8wMsMFXHWYLfDvlazFOG0v8m2MCHHDP190njO9rXjEOjm2sIQsD3DXMibEcwX3G99zNxpHDN/g8xOfGAs3HzOIag+PjeEMuAz5PYWPFPJzAxmhjMNhY4NvG6ww43H07NRsLfM64zpzAWDCW1ed2ajZW+DyErGoc7nOz+OyA2QLJH1zj/PFZc9ZaSHYaxzzENfT6WIF5KBnC2zQt10prkmsTyhXrMBbKc+b84Q5bQr8wllgPyjhlOEbow1hChyW/tga1lh4zpAzh0+GwOeP7YznyeTixsR5jcq00LthIGdqyxKXGEuuxHMV+cC9d87nXZ+krx+LzkPKUfqQMxwLsZGkcyxHcT7kXkTKibpmNxeEzZjm3/Ezs0ZOQwVi5T/hd7R3fuPwTZoZ5/vPvWud6ydU4uuKSEOTgxohJui5uSyzaWECtgUvpMeMeUn4t+jzAMWoTc/KwAedkcXQCW8/BDxdTabAcyQxQ+bd2zVnX0UY/uhR+uBgGaQzpG4e2UdEN2E4AW+L3vH5ocI7HJ1wGUQKcMw2BreeoBDPGsqyYh4vwsaJujLgGv1P/pvGD0fgNYG7aRnFdW+DbyU6xfTvAljBSPgawbfFdKeA8AOOIMqlrYayweQiF2i5yMxuVdoH5lgbG1nPwuTXD5/zobPICsB247iijqk3d14xG2w8naeSldLABl9JzvX07TV0DDbCNNfUwlofKzM/bssZ1djIcwBhxXzkOG5iHixjruaZWzjFY6irSODlMG3I5gm2noZMyPDToYzmmsQ/9Me2Nyc/HKocRyM1OA0Bds+UoDO1yFPoEz7mkDOXwcn055sF9lLJHGfaxwMcpnXWTIY01xkqZHAO20Ngb1z3Wx+dp3csMw/3qNd60FIS8QHjENSzMWIHtNCYL502XtCvGxbSxwEyebJTHtRGfl+OXQthCr25EH0irG+iFSi8lSlsmlEMV1Wa18DSWQh01XowzCKdZ0PSQRAu6ri1w4+abYTRBVOU556MwdFwQy8210GhJtgb3jZ6jFMLSosvjLtzMh9h3y3FuFrMBLLVGxjnGxproP2l8fcYYeb8YklGvLL2SvLSNJQySFDaRhTXPV+sY8vS6J1Geo80JK2CHQkfuJUMbidgS2XGdgAnP8XE+8ro0up5zkJHiOo0Fxg02luNco0BRs21g4zquHLuXUtsC2JbosxDurPt7IW7jNUNPvMbk2nPt85SjpZ5Ofpy61KXMDe66b3N4bkNmKTa+ZDhWyjDG4L7VnrFm3DQGG9QRS10B2vqPgRUAzGV2PG8Qc40Na4SCxo3veo0QzyQQD6RhzVPHglBohNCwAfOJOQ/APA6ryg0MF4zURp9xP3kRTcY9rO02atHlyWnozL2ExLAhPL6Eq7nzRybaJ8ytILestwQHwHQ9/o68NpXGXD4nEYdJpmMBMOB+KIWzpny+RzuYgs9IOJubJ/80uG4W3nVOYFjJzSRPridAuXNzu8MPp4ksNL/0fvyO5uWUmcljpUwM2A78bcCh8M6Bybmaxe+OnKvW1eCFSHNtnddjSLkI5QJmnoggjQIW6mnoQ8hHHjZ9cbwuGSrkgVNHTolsLdCRxiijJbQ0t7quTxrbmToRRnQCxjl4k6F7k5vCNXr4uVHPRjkaRyJsE+JIlI+8fq5vXkcKTpnPSXtlec9Y60DQfnoaIV1eD1hTSIkYCJ3mAcCSe8h7zLadEq7PUMqlwXAurGJNn1sqiixmxtjbAT5O4m8c4uaL7l+QT94kYtuVCr7REyzAdohx20jrXvdz+OEMB6ENMuU1VgBbvG4UGiGmruPyul4L6ttpbL6MaAjbp3EOG9xmfi+svkDulhtXUDW/M2k45dH13eWIMax4lZnxuW9S7IUhzSDCO861S15mWWm4KWvBWSp7hp2pYIAfTnhvT51ITmFyQyg0lNy2Q1PE+Letx8BkGOAe929GuDb0LO4rwxN6/Y0hbgvl5HWdhtPnRaI53lv3ov4Yjks/5gbbDsURACkD3w7ACs7FgTEjDFpH8gw5f+NayoHSsDidoW+8zqB8yK+UjORwZhqy+O5JGBcz+LZx3t2hEAlKLym/1FHO34wywhahH9G+IgHZgck1DRkOrvGGVdY5dMlCPxUaAEW4LEcJF20chcK5Yy6eMFuEGWQth2DhYFx2qHDHTwmVVthyLpUyyKGR988xJJxfgClYTLgloZG30EKntR4d2np9F+ExguQbwGZpjFxEEI1d+P1BL+OBCkgOJY8RgyiYJ4/I6wxbaPoXboBOVoWnCBCx0BtzbcwBX2CDsTA5DOAAcU1jOYaPCnNsOcI8CJIzJCDfM8ZRKVqGAUKOMe5hR83I6D/WDKZz/RY4IkQdVuElxpbEp4NOYuF4iDR9mxG2+imVVWEBl2ksgRB0Td8y5BSUD4QBhhwxvpmkctNHIAzpskZIOY4SpcDI4wzLtXF3jPUcpl+A2YrkEMmp2bJiyJCal14zpInQYQk+zgaRisX3OZf493GRtqmfRA1DBGiFv1h4nSSJDy0UDJ3IMFMoV3quNaS+mPbEOIal4Qp9nX5aBm+swFiwBkSZGd/K+06xpX1Q3AhBhpHV9W2XdYBzQ8wJnxLmkpDSc59q0217y5hIh9DKiXO9eAxXeEJkkUwyPO4pcjCtNC27tFBEqd6fDK98a96S2YwtkI1vh1AOLnTLfqBY/UNbmEHitTzmnBO2HkWYYUaCMcbkh42v0Xv7DEKzkbQ+iQDkXUJgJUeGHS7ysKEgYnzIk3qH0KD3MAuuxMJLxlclHyPZK5juJNk2QuGtvNCYiU6dPEaitMmxuzya0Ju8tGJ9Zg9ksJbjRF6BMg6Nx2hoT+hAofNYA51mVmkLL6sMUX5buuhwt0JdXmtUYSz2MhQxajPHEJyJM0QVslVIOmvMuvdWGSvxfIFsqH8iRlP2zOBth9CTHlpBexJItKWsi0/Am66Cc9EW9C3nBlIBZmHMVgO9tlAARnCBs0FuerjUOeldwiKl28RyA0nkaDHJthuM8ZvVRp2TizNLhozhA0rR+rvHRmLYoYkGkgEhP5WaG7QMIJJ8ihhWlnbsP9PjPweKNCqr3FNiRq8Sdp1enanIyop4fjcNVaqpVaimz8hLzFkyZawamQIrozg9QjiFEVQuuOQr+VC2PoMk9Y0vOUNOKzmkASrjkiSyQi2AmZmVMuzKSrkmp6AwdCM3s9APiHG3WDdd273Q1TjKTRtr0OL3roviCDBgkB4J8cnxENYnorBcH9+I0uDpWJJvmhvlTP1liYCcX+4F8RhjTR1URimyWkdnxsrNKVQyt0IINshtIOTRHHVs0KWFtNhlKgFwvUJ3xnKEebhY12nRxO4nObfSAcASGa4+T0nI8LYDjIWZnnKEdXR656nJAMrFwj3i6e2UsPJQCkpvlgqfXmDy2rOuwevm5oc2ZWyiuQlyBYGFRBpnJtzuoWvHa+N2ynP2e4lGuFkCHnKRMjtQ33HfQkmSYLVERyGP4isSKckzTKEmhmCj1x6cppwL9kesqs97R2Sag9h+zltxeUDyFdgmMAKBZSamhXwR9fhuI3WPiiT0KnsWxk5K5UUa0jjJ+zvJZYVuAGITnp0HAHm4jnaDaD0udAE0R+OwYfJrhOIb0Mj7/JkedFymxVHIa7dOoYPWeQQJSWiiGX2RufEdpHzC+AlV8GZeMjQiLrT5wA17PmmWAwDgG1FuIrYzBl97Q/rpQbgDDvOz4YvXdzV3Gqx06ADWMY6B9RiClUZP56vibnnLc1DcLyKre0fFzoKzdWMtRElaqbbclIptfYPNSvOEgRCpqShb957cR1KoJbMSnoQbcpP49IipEYshNAAg+QXzAaX/sCBSv8q/24AtKwVMI9dTqm3jaS5DMb4t9XkhLjM403IY8jK9IKZSpCU6bWxPo6ONqjw9fHJ9ttzoczvFLr2ahnzUOsQil4xpTKooagDYELtMOkEjqcIuzW85imuYhQyXIxKx2PFPc2PqfColq/lRhmMr1GX0lkOcDPkSY6gwLDmegvLFf5QMu35KnzZGBtzo/FzqFoBesGcp/+Z4IDTrpe7NCEaY4m0NhYy4Kc0TvcLEncU4bKzlEmXcxM1N6W6MJWpl1kSDFYqrvCAQ31gviT02jsIxZejeHBcNptY1kMXhJC60Ib8QsAlwjxTK3E6DGKtKyhC02Nyx7G3CnDBT/B9CMSCUsClFewemIi63TPWY8r8yMNuGMYqtNwhpNITChTQtkrx58ixCH0IChIoJwxHFUYwJ03LnpqGRktW3pngAFLoUMy5GfGZ+Pxhtfq9V18VGkV5I4YXKlHKcCVM7XDXG2oNGOpXXVODkbW246bwhGgeQc+H9vGQYf5cnz83tkdXZVS36jDQsxLswBCAJ7fKuMzgrlxfT36rx8XComWYUsnEHxtyFUE59USoaXH9A6UIWuAl+7BDA3q+J1A5vHnomtJGbGMCOTFfo1orZMq0+RdIiw7Go6+GdFTrrZ9BQbQdgYTYMSONtyxrhJ5DIrXhAZkGWLdGP6okUZvjhFFhWAtHgdDKkH62aGbHW5o41y3S95ahtpNKE9SFZI8JTsBuW2YG8sCzTcpybHbZgjKPwcMyiiDAzW4LhpRIChpH3GWSoGf9CJM0WGwAqstmC3Ray0dZ1eb+wwkF26RqOQf4ivV2HcBYxX7L3HFdX2LFwTj0MoQdX3BrKwJSuaj5yTFSohajKKv0IAGORUQyySfF7ZEWo5IyfTVAVQi8rjdIKkcJjrJEpyEyQh0fDSLRVRUHczGNBMvm2pozHUIHRaMggrE8VeNGAjCX4SlWexm4M+SxrRk25zuOooRyOJfkh1k+oeI3hQyLTHoYBMU6AsjhCZriUYvbaUIk25WyYSRpjTRsxxoqpwivqxY5vGqyCpRFwhs4YM1H5GCP00CSKJd4nUve2fkH9qPAKTc7iiXyPGk3IQPrrtCMMWcYCGwM2JoayWRZjs2UUkiOXCXeMYcBYAwuZKd0YQk94KQG4BinbJwgmTyqPAgrdGoEoCz/zWqmo3VPyskVctfsJ3mdYVDCynwkpJS9Pn1kCxY4N/6QXjCuR/Cqvgx6PJvFmKa+6P1+TobClDIjQEhSmlXdKPoH3kPfQddPwSSbyYJDjykAKWdyzWzvJ2QtlWYWWff3KE3eUtEcKcHk4XRe5sbpnSw8MrfXMdePI4n+tohBU0Ezj5iZsBqZBYsltX+1oOdeSobf7Y6c3pS+gDgNZaIX+R1dvpegdR1PvJccM3VKPnGJS2L2lvHNM3difkW+GP9bHon3bwxlWto4151ufaTqhsWt8uzVr93DNOcYxBE0yVkvjQEZ/znZjsfhkY7kRcqNoQ/M6dT0aIaEUZTogm8GJZF2GQpriAwRDs+Yhx1ITT8EwT222ZD5ZY47LaqOPHBfgyUnALOef4xS0VEZjFw+XseyhSsqwIa/kR3Ksbc5Zx8JaAtQiQyHHWKEK0IDGoCLps2OnIFVCztfSIezvX0oo+Vt+x8bxfn0NULl/R225BvzM7TI8SZzJCKNsZQkTWbGqDSi0lAh4zfmHjNt9EnGMlEVuZgBCeUavmgTl7Qxtl2PpoghrzdNSb0sP6j2kcR6sUypHkyaTeyU+ozWrQ4ulq7swqG94GZbuXFuGDTmv+u5e96QLGs+S+y4RsMPXHo9HnbnyrIcSlAUzOwF9ETBgNs8sGKjMgOvQGN+fB8JaxaSwuq/y4DDANkylpoybFICPJdI/5EhkvafGPxb4JEELT+gpRJNWu+XOk5fwVmXJnLizACjjOHhCx6zDYEg0EPAtdZ5VmFmLYqxHQDM6w9u1tfYdFfUNVdWfm2Ct4tOptKm8GVOUOA0egWhHHtEPJ0yvIlGBD52nAdN4hOTK6vRounMvAHCoSlfNwbcD+QqHjagLSdTkzGyA8xeHswQJHelUyTAQi9MA+zxtZzqIPJXR0I+dlSEgBKKMg88Dq0BRsushLOdu3AdjOaZux2HEkOEJjWMhQIVwk7oWMjxAPIU2bJC6He2Qm8m9NKLCcmvEY0PHKQOQi6DehAwn3Fn5OrV21F0gdAIgF1drOtF0URyaNnrI1NbwZEelmIwNkR4aMFthOKSn1BqMJWKvOl671gBsjdgo46oFrrpoi7hpnnohERiCk5AlpWVbkDAyDgQxPuP5ABsri77ofZY49GbLUTDlTEXZpG9RvQAQ5a5mSc46Y18MAJu8TfAI1ja+wYiOVxrM5gkU6wbuL8tMBVDFoTxVOghdfxyhV9vRLSbSGsrVj0GJobxERzA2alwOmPiHlbKVAbEj5CnXGAjXastNInIT5KC8IcO+AeIjJG95UjPRTSxkeN4lzu1goFWTMiOgasWxAlJ6tUlg3J1l/UJbMp7aUJJhD1+APE9iI+YcKeKl0veouUTUuFTdhI+c/xwTxiIxAxJ1wUZeS0cazNaoa9EBO/fSQ/FflGNlIHjPgSzKSuOTBoNVoi7kyeyWqVraUpagM/QW5u9QE6MAG0ajKpmXDsMGVsxDWMoccFR3RX0BBT5VYaaYMKzNPGy5SL0aEcbqxbXOJYz1XKINw8A8zHyvyooZq80ZG3Zwg2nSzExMVpP63JheO9TGo0eH19kCiENRilgjpYc0V9oLcByIEsTuT84v0qnGYp5EBTq2rbE3yJ3H3NvZEMkoz1/keYXJjEDJQmST2O6oMYjPmxsmPR90ZoReJ+ZMeWwHqI7BCE8dLSVoFmd9eijDI+WRlmShkBRb/FD+N60der2EioDq/a3I5cwG8T5aIyElyRBeCGAn34lKDapyVVm6pWSY6Czguw7EBUG7poxVTl5nPfr5nNDTHX/kG3y7iOrXUSeKE6WqwMpnHDuaG4/3OzIc5rjqJOtR6QwAP1wsOWeUu8WsWGG5O8OjsfE1n+FoOqqScQ3UAmTJu1MXePbID4cmPwCHE6xwRx4oVvxDIiaG3EhDFYz0nyQnVVmGtNgQoZjWv7PpCyYnLsscUHVEzjy5j6UQzYiFGG3Dhx4tqUQgYx4FMhUTuvVS8VB8a0oub6uNis2jWjQhGWXA9FfIQ7G0ZXhhzDAk6eeOPMvSSreBybLvgTxZ2QplkrhNtEBZ5tFjq0yUI3mOnXfU3xNQ9SMsMkkqbU4Zijzm+u8bHYmHUe1FMx4Jkw8VV6eROyUqoXdL5CWDWpW2hmqC041HGg2hj+zrUEZZBjVhP3VBqKraJIhjOyqvOkLFSw/r9eQWxhpOAjTGc2NmSXKNL4gLouDq976PwDXLUnXwlDF4UpfypSGyXoFLPOc+45xR5ytmVfbG1pv79WzhblU9b1BYmE5pl5xgtivAM4aRgU4yCoIoAdeK9d8TkyJBiyRqCs0NoY0KwdgW/2ZZq9Dv5HH4Toble4zL50w+Jaw5uQ9NXNBeG0DQUK87duMPksyQRGJ+fjQlKMJvz4Jr0yO+Q8IMkiLvO9jvAtzQOxnys0pvlqEQKSdlbCHJnBSNl6LQWAndiT0vObJk3uO8TiJHSNliHeIznobHUiM6oy4CvP7unwPnUdkMS/0JUVVGy6CUIOWlAjY0eE2yL1LZaGvQCMJ8nY6Ca4uUR1t7RyKglKE4EWV9NJ8uP9epXOrxdqh6j9TV4qFyX7gkiQyXsi9K1zGuI5rcdmGv1zzGOEqjZqZ6m3LKSnHn+02+Wpd+jySQU7ZtvVWxDcOaZI+LTOLm3tpx3ZabjiO2vJiKmRKO0RMZDwDpWLmNhHbJPosElfHlhBMymQyHvH1T7LSCCCPBA0vR12DL8RRBx5/Be8tbCfrDc476yVOAJGDj6HOLgZNUnCzUK8ibMHDb8jrVwCegYmZKGLEXTOzhh4xiMdv9yH8s5pYGJtawnUchb6G5hnF0KIeeZ3V2KGPkvz1RQRQxBzKrEBBoX4NT/hPOsuQKXWOD7hCDvkxCstCKQrUtdcQzO4LGr0zMedo29gYdDwh9U3imwqWeYvU8Iq9x5IEt9WNxB6DQiSixk5KgIe9zUZn7kCML3YkQR5XGvEfbS55oqXEn1nSMiD1koc+2g2ltnaTbrjJ47lPVkwSnoXqjUW0A+jkup1YSSccBvom1LBKtl05PEm1ESLXmNMZ6nKjARovRJHwu6hhHLM2lhVO6qx2uGkNdoGqv9SKq7sHKi9GDkQyPax/VHPinHLJiSsalcA7R4SomMlrtLLueUYTCIi6HwRbBTOOacNNABJ5QFFIucQKXKeRuOPM6qiewHXgI3eAc6YFdoYapniM2DER4Gr8jr2qFSrIrlZc8OupLD2d9LmXIAiWmsJHez72MeOpQOBKVmMvj+wSP6C8ZPiVvQhlU9qYZB3Mey6YugGFeypBGcNBASI+GWh0w5WuxYUTm2zhqmR0qIDez1tggnSD6pH7skLSKBCmzbLGAIPwne0goLcrBxefV9i4P0e0Nkc5C9Ron03WYfCgjYdRv7l00gncIqVGGxnB0UJcUQo4gYnNvCe35BixHEYbkZkyrTUVK784ZOGNzWbN+hLfHT6jPZ1ekHVyjQuq1hDqSlCAkw5c8pXnmT0JojWemJ83j8Ypr49Ua52xjdSTqqfwzoJOdYVvoOQTjCAuNCwdBRbH0XnA8eY4uJ8o8Gq6I32jvQXKieiplLT6pGVF5g/qcYtCY564YSwY45Yg2Nsqwrw2kkH3cNRmRYyEvIbOWoUgCro7Om/cQRUz8mvc1hYIJmdvnpT87GW4ZQtWc6r4lwyXHaV1Vc276vgxVI6udVhz7UGE/HtvJ0PvctW9yuWbJTcfTG2JLPbNqdF1R00yEqBA6wtng6rSf9jUiFY6k05he85tCgp6GpfZszGuNfGw7FUhiEjonDwtLPiewcPMMHfOeRdTQOprzHL4IF9+aQKvHRSqXcvpsw5bQVwqUbDzKm89TJKmFyASMRWmlWXn4uXHZtWEURsRCmXSpK38SP/HWlDEU+5ynKUH+ZE8UJjkoY8pFFDzsCMzgLL9GbXrChB1s1aKNGGuGeO7oDUsynCB8dSKksEOtWQ948rOFlyIEvX2/w1qNK3cZ1zHDShlgc0Q/C45/WcqDpw5uaXjT4ACx6c0BKxToPBFdDYFUo9CN9IRKr6sGo2WslGnxDWaTXvsEeUpUPAMbIrtJ59gdTFqkUPxwAqwMtRcgu8vLEshIQhsb+e9iVCN02jmClOOMUKY7MNfZGu4jc8SZDu2rrcYo5Ky5K5s3liBRVefRUFNleyL0ixJ3rU0Y+XVkpVavLx/pzXdVbbKwXgeKkhDKOCeUzQRhqVtG6xVt0znpsho82+AYC61whisoCMwNWEfmdS+gDokdar2o6Eqr6nCa6++5YdhxKRSQp/e0QYYVO5+5Z2t9JWH7TSe4KAiMSjXHPFt8yTtVHQPytTQQaOQXDZmNY2Ycmgec8jbcmG67a0cCpvVjoEc2nyrWaJu2SqarBN1gCh/aexmCSOiIMQ6RtUKGMi69ChjODb/F2aHMwsQdh41oPeeA+mAUMV5rH3UwHKsB2ZSG76UO8r++bRir2ush51BNfkKfxI/kZ6SrzFzFxlYqc4MtYayMPTszBE0dVTZJXBE3SNsPQw5tlgwTSWZ4oKQCZ5Uy5NmfrCgNPXQD64uqCjYM64QNphwSjfK+Tb+km4EsPCrnKn3ICWhCig0JR/KAZ7pYVVHynPwYcO8k2AbzSilR9TCVKuVmHUNlyWyS0irV6B55EI15di6Erp+eR0eOZV2zM1GDV2nMWJwUlVgQfFSVZn7ea+zAvgFqepGsek18GdfTBqbgY8GUD3eoga4UVDGwp4cSsmhp2yRlvEIqMe30mPHSguyZoRBlLGyAU0aqjB1STt2owSK0EzrbVU36lDQT6mbHqkzF6aeRePwuhGo1jryHKhe5Worrp+optHZCsCRXIRPdZVTEaRrV9OiAEKyxYLAaOYsL6PMN2DnYYk+1D7vsiAy5kE6GdK060gu1hHrTOdJBV62H7eXdUMneeDdkws8FOqjHCLiru1w9syVrRLKSW0iSBxs5xrVzDq7qO6GAIQKs0qfR/qxiuWzUwjhTGYdeklwpIHmWGMBQ5WiCDEIiKL3UlBtG3o6koio5bdAzjrDK8uA8GDdGt46m/9MIKp3Ha9EwZroQZw3eKkGFkg5LewGy8N6Of5c3KteWR5opr2gPV3GpOpcBYM0GSkZmfDSBKlY5hwbSco7VvzA8KIlVqA8EN5yxp2OSXFCczKyWIQ1goZ99mlfkMYQOuR2rY7mMNaCYWa8V90KkYGshg8w2OFpXZG5ejaRI9hieTgxzLYUa2rHryHhIzl56AGYeukBThkR5Y4kKUYYG8W/LudugbkLrtVSoDkc+tsCROlpNiKJxVIXMRPTKHHY0gbMGu/QQO1Sn92f7fq8BsXTYZRQ9dSzemwCGrzt2G5rAlpssFHyt52SkMoWFMpaYpn3L/VHQMIS05ARkQffVekAW5GgzyjPQkFUadubmynZ7uu50roXT4422GGEt1RhGyhAGaOyMljxKcjHKRMCiwMsHMmtjKvPlMWox5OOoFskYqwJlKDBLhpB3bt6CxqKnsKUkyQ3x6VypgIv4EhozFEI0cgWeSFFhRDN66KcfA2Y7jXSmsoVqfAKo+pheBRoZGDqJIaPIxwlIFtqrg3rX6zSSyV+5thVOqugrZFiHC2OT1P5JLw+gvHTXU0c/BxXZKRqMNBmIZAEAACAASURBVFK6BoH/VPUodXtWaC69B6qaE0ARh+Tn5uwcB+r6MhBJ6FZ4krrUnKS4iZgL1yCziO30uBkCGepo/gI9eErOt/YCam9JF7U9rStnQurUHG4gKUR3Ybb7XMVQRBz8Pb/TX0sIj7zfLmMCK4PgMgzgJihIGxnHvrnKC2qTBDooC0ybh86yV29Ia/PgwifZ146PQ5C7hTN5ccpQVl5QBl0h2mebAlfHb+wNRm7UvWxTCBnX6nehRcpO+X9QwVusHvNuY8nN3EIbNOOS49TfBZm7t9pttDNjSIieaqf1OauH2N8zOTVV97b78Hs7kNVkmXUuaPJrSKnaFUgH6ppVFHgoOWV2o+Rn+5vv9oCl02sGOu9FGbbDZiVGyZC1KByDWWLsGCN1uK7djxfMJgONiQ6m3S/HixYRNNkmZwE/hDdO78UycAc8T6QRbs2tyCAuhkgmtZJ3NbaR5SdEj1GNajsvqJ3IZgC71ur7WE2twnZmS54Fus7YLXiVKO+Vq7pooRaqwzVBS20WFUuJoyGkBZnq6DMSLHOuM84YDqKAsJEz5Ry3I5Pd044wijkgcKQIKQtBaIVjNOgVCDSPlFzRwK7eJDdIyG3X0MVJflk3olFSrJ/ke6zxC2zTZpQhFAok/8K5yfPCq8+ljJrIQa0DzzngIKMkp9KLkzgeyieNiYw7kY7K0EWiJ0dSMAd6/J25x2G3djBNaNrodGINpb8yH/w+ykCKCsjsB9FLfF9P+CMSVANhZTtKK7m3lKIVsonXQ4Z93kIIOgPjmC6kM2A2sXtQUR/X1Pfj+mtn9A29zl6nLT3CEPRmuUWgpbIJnsrL0QCl10GvPZ98vYgX6PpQZeeagtJE8gSeO9zPxnCMCWl99ZCdiq0NCfUp3DxEA5TnRnnHRBDqOiVoB5bGmpEIo/KMeM5FdW0qD70v5W6hAUAvRSUTV9Dz8lISfjaOu1NRdrFsyL4TYx2Ki3jsZCuM9x8LjF3XvTURBo1T8hLqxGRLEJ5EAXWWhHM1oaA4nj86xIZxU9KZUKeyP0UilNiY8VyOmlIYz1YrIqTq4HrQEZ091wMAxtAByqr18LYOVPUj4RMX6/pZcSnEOHIdMvU8AOi5L7OHdYAp9WyHdKDxzoYIkZEIIHGL+BEZq9Hqe8ziKH0LB3utkBpRuThFgF3OlK2xVs0qFMO75xmn+HceJJOFDm7gsPPMIbi2ALL6TqFI8dwrW5EL2eC7vpcdknoM3M5jmJquDLgLlWzQQ21iIfTk8kIPSK9JBEBFKZNitbg6ian4HbLeIvK4qOwPEL8fIibcvTfZ/s7LCO5kKMNQcWDwGfuQR6njuHbNM+S/lWcyLXh79mdeZElkpg2cTVu1niTcQvmawXBPTiSJLvf2LNEmySRwW5iV40cgh03eCjTuKlMHAd6ZjAZrSEo55Q0lk172Ln7kTNiRyGXCsOb147vy0siwoBvu2sxD8CDeG4PIYqaoTZXIlGeeeka79hnjqX/s0t2QKgkFNLSV8670qZscyaHK3v+7ZHrJ0Oeh1oUyqn6nDucZGju7ppJh5mtHZEN0fiGfh+Bs4LGLEwdwOEGdGyjWNONZGwBO6N1oaWWIoMzCUVgzxn1Zzw+E9WuDdpdVJBHVFa6Pw6ScAzAefU+iVBvdgSHFCbjr8DzBqhMkJdh2fiCfWRL5bCmdFD0fFSjFYU47C7q8vu8b2wFw7p5PCPNSOj/hWLam8IjGwCRONa/OiAdKKcXZpX/hbd6pxcij4zbqeLTkpjmOkL3n81/p+aiIyla5PNNsD2FSOpaGBzCYCZrH2js9X/JRWjMdPUglBhwzyXbV5eqxjekdAbhfhNKBqaO8AmDst3GgXDzIX1fhky5DWdyOHFVYJC5iNmQxoXgjwtXTROn7sMNqjbR3lMps3EPqby6y+oTONPByTilDC1TvQsCzzs2gofCcn3i5/x7CkG5vJ/H4wnwkW8KXQhr5OpVisrFMNgyxOEar9vV59kPoADQCfPSeHlUfUHWm0DrklifMgiItlCOtrCbSSTZBMz3ZHPMUOgvQq0V1NHwkFLZobqNeHjkQwPSEL8khNWlGWszjtZHnU5jW1OK45xh6KjOO6wPZn2Kqy1h5fp2zkEyCs6AMRfwJpmqBK7AFfACDmSVTsxyFiKEU1T5NG1myZNv97STkieKKvMlC6epEfzL2ioNvR5g2GXIdQu1W2JChtZyLsVluIoiU4ax7jcnCL6FAnhWRhNSzxAtJqglvOKqGlrVR+V4Qoj07B2QDm0Q7EZ5Vy732iEXqdhZbMTQp4n+WXtqAjz0qyHNGIpoRjBSaTINDYavAqQdCeUsbU15j5RzLAWU1dsqzjGNve2Bj9dXn1p5ixVAjhROTy5ZwLq9dnitTRGndC5HsC20ihPHDSaEBKS3RQsJh8QaCcIrZgGx7nwrFBR2tAUw+sLi1HMvPs4zW5ymyXiP318zxV9HKGaTRMw6aO4yboxFvihVj52gygGorrMlmEAXNQyj+WRk2qOqTD7VtnoEQIP/KVLAWmkYsakXQDIqyHJyPQhsbqIf3bDDbUpbeNpRvJ6G6NqqxS0J6r5Jyb2Qdzq49w7btsD/f4Q496xMOzHwSu8JlQWc6lN6+DgB8zY3pAPKsEVGhox4HqM0fRx8KOckRUoqJUHroI/I79gDHkIRhe7Rnspsijmlg2doR5Ov6po1hC03P7MzuXKtae+nFoYjRUK76HPdJXFvhHVjBqzKE2H+JwnZgyiMT31/Mf+Si8QJzIuv5pVziKXbxDr87Pb8bAiyLmdmL3If0wG0ZMqXUCkakiL2wK3RX5cSV1MypkDzMsERnFs7EcfmH/65UnaByP7rcfmZ5W/Q5qZdCl+xkGNHnnR63IazdHxrpFvpRdUtG/fNtjD2VmUbtTB4+uSllpnRdhVpQ+Njuk2ntLkONQXF1M9RyLruK2GZYRCbuMcRuXioccoYtJcOONNu667Uz8L82g7X/jd21DMpceMoreRLJML/XrtP0Mnt1yHjnmaLaO/la6mjb5GjkJ/dT0Ch6Too+3xBKTl4/7XMpQ11va927m7M5q1O6PybWMAJiZvl4OMWbTTkVP3vGzApDjGfit1TC8oiyZNpwrQkuyoJZgz/G68XzDYBeHTi3EyyCm/OALGwinE0BZXFWeMl6FKBh2IqZnqCVIXeURMXuncqjsm7JcUIQ3pVKPpBTmFDx0a60F4A3edgEdnwOvGS4jB2fU0iFY15a2kyVlxn6hNcIQngk8ZY8w3Yx1zgf4oPuLVt5umLuhS0RiQR2PTydGGes2DVpFm8xVElbvVMzDtba+8w1LQRC2C2Es7W2dQBbwCnGlmyRhizb9vmEOKcMlSDjMZteLimBMmrFB6Wuw+DbSYxbIap0ACiDAgWv4i3UAjBeM1Y6Z7k6H0QezaqVyXHMlqauFK/Oo6hymht+6mBjG/JA7cdWBOm+ITrB6f2aY290nY5mTqxjLNF81D0a4NqIODLJkJjQ4INf8vmdaH7c4sEvir3iNauJqD5hLBi2Ru/T9FiEXSZvN6DwQ2W9uv6yHMfBLh6aCWspZl9lz4YBGTTG08tx8zyOgZFNfhOxZH0BjaP1IiNE7YSxYnCpuo4IZRbCcOTYg4/pbPyGoYfsZC9SZ1pQv+tsjLIPM+te0usvRyEDnhhsqhT/Z1waMFdesKG/cZxKEJ/TuRhu0CGFjJcWWIaC3rXQ1Z+i3s/+GdShKlv2fL1keASVPk8ANhYsy7mchzxmPmhpkddWNycZ0eJknKGLieuxsBPoPJq4K9RDo5S5M+ogf0mDNrLZLdc4Ob4FqkXSd6cMI1fHm4zcQ74MQkIndjJktYWyMe2nh125r5bj1EOkDI/TIGQKVvt5x8esueei31V8XieVzT0NqAHAWIPgjImXVzXpJuhJMnWmcxvKEjBFRJ5ApeDUylzQ7G2YA9ZkBiJuLiVMhRRxmbXpFD8hmnFsTqioVGlYfD3Rqk4wZjrJjWSY5fizg5eO7ua9M7iAq5YiuyVJQ7zCIIuaAgAwl9eR/hdkVdanlIwNYqhEeaBvHCf6sXEEx4RvFWIknNZGSSiZbiI/tz+iX/Lth4oUemQ3bX1OBjzRoJVxTgdB6s3aCV9r44CIYitPaIi1g46kn62LqdCheC2tTe/Izt4X4qNQaFTNgRxOR2XN+y/IU8rLSn6B8skwxqhvTYY1rUTTyiZUCpVGtz3DNPuqsklPNNcZZz6Ptk7ScR0LaDpF5AQLMtfmhmErNo+HTienBSRKrL2gSS65L6V3YU+IztBKHCwo7oB4uvmwtkCKObWVW0mpbj3bczxhLHjxWIREJnz2wraxY3TFkNmt2D0ONTmCwJsbLb9qNgLOwY9SkKoFsLGyq1AUFMWiE3EsCnss1dY3ppV85OvVl8Khtu8yUq6UqLweU1EqulHdPRiGZNdl/bT4T5Wieop53LJSjcjmJWBKm3M9XIQKgnzTxiYEViw+D7AjwkySj2O0vqcwQldlbFChpuCxLYxCDzneYedapSSoaNVV3fVYwe0U8Zg+Pdy55q/cfiAuZXgcprQ0Q6x6bqyOo3eejOsjjsGQHho2oOeTQOsCqzDNgbmdQEjZaVySq5p61stMZJDd57V23Di9OLBguwM4UJ9HhqRgdk0FWxkt8nch9ZRhR9uYqYv71GbXqy2dQRL8u1OmZ/QQ3alMRCsDHmTkNbw36aaO2HS0VAAnIIiXg6q8sEN9A6X07Uize8RSer5CH6j3gbafJIwMIz1YCC2bCGdMNsuLEyImc+2O3XM0c9wqZVdI1SyritAaf6L7RC/J8uA6eJZWnSRZFTzJeKr8W1Dv9jIMZQvDNmUwsqmJ5EpPKUXN6+lWWg9ACM0NCe3zgFoefstZR1sAGxUfJ4LgJ1IhtZE8i8+CIOPG9DI2iRR8Ur+r9LtkqGvo2HM3CqUnClOyUjiVGkRe2kTOQ8kyTrPkwjR0ooAI8JuBxc6Aa62yLUJDx0OFbWDKEoUEVazlrGuwzCKVxGseXS+6Ptpehi2rWLoIrrbQTVWYVvFj6ZqMaWb0RNAnupczdPhWmU/XKW/urzyEmdJoRIZxIsmQS9JdeXYbvsqoBS/LUBTzHWul1mHIzdeVcaoMOUmnQ1l874STB4yTBRZZ064npGMSWHIA/adZWY3daq79UJfiyTI3BekrBOg38JKhFKP9naqUEFP3dd5HiKx6dgDyGDG+bEYs8spZXJcy9J0MM5Tr18rSbyoplTXGU3LXM1SaVeG4PP/mhArWWshQ8oI2L+hdmzTPzj83svG7/ffd2hWyONupqsK0WXPUdWk4tIHlmeVZQcLaKKeUr4scnbk+gXaLFI+Tz9tOz3cOZKd/2I9NusY9l1g49aoogOr6TkkqnS3+zvf3sH7PLouuh/me7tV02CdGlpPqthrs7RYTNQj3Si25Qb0GQoF77r4Y/pAxYY4UMxdKyk1IpY2g8xGT3k21+/R02f5eYyGUleWVx5r9eQyy3kRS8d0aby6gqhWlf4jYNeSghrla1OaxziKYlCEXGURjrf9hyJD3EJTk9aJ1/2RooszBVrLR+Gcpu2SoRyfofi647MjfU94NSYTRsZSpOTC3ffpUBrlKvJvHhtW6oM3NEfPPHpxAD7u6rBPxNJ20NLZL3YP3DltDec96Mjpyvn2epSu9zmSvh6WbmaVJ2Xi7RtNprStQB/6kvzJE2rMcU+mN5uElw5Qp9j82oMOSyb1kqr5ClTIaY7+v9Vpbz7i9t9dbjQ91b03Po0MjO8Wh58x2Y+wjYB1WVS44y285SSNDHpVoRwArNqOiEXWykFYw8916aG3Wv1NJWgWaMe6HvJGQARxx8FP9M4AO9ZBerQMBzpd5bfVJCNJycs1b+/5sqSbFmVwsevAw9a1+QPBUBKilJ9Qx/Ao5ZKBCjgGN+0nb2ChDD5HmASIRfXltqwdRxxAEMYWIljRg2f6+oaXoxLRArfmrdgLJW3rf1IamD00RQZSi0u4B8huMq41oaaqWRVwJ04spw4Ycdn1BeJsdzDfosZnSrZHPrUWTUxDlM6svi09RFgkGNmlC3b+jgMX4TNFGkru8teSt7FnN5wzmyilm2DxaKApAz9lNy9GeRpaH07pBQjiaqF4Vp2all/y99nLpXOw3O9NKYsNa0JyWUuSKeyi3UIBOIpLQS2UwLpSW02ndVLWYN+d3BxCxly55QHY2YkjkeQ+0TW5574CHKsOVysr8NqXyyYVCGbw8Hu1cNE1FLH3rn9GuFjqqeYqcrUXKIi4pKV+XkY3PoLxhhkYyDlQiobg8Li65yBCrYxc4/s63eK6Bkz/IoSAU2Pr4Ukb9PgVhDbpOQdQ8kKX5tV6kOwJOYQ83Za6OA2ikNkBDu2A/B41HtxGUN5JxJj2jbU6RV8pQhlM8RnEnmrelsc6NzGfRWvespue3tHXm56v9AVLHLa8hUbYwXShGIdoZGWYJQg+P4NWPU05hztTDdEYNTe2QdEKZGovAAIZ0oqvb7VtAAIbVYJ5dkgeSYKozDuW1YtMWaztIoLmUi3FqM+iAxVkM1a8LBkUK0WCo50QUKeqQB40Jqe2cNn2fiOmX5oAM6rEQ8wnBdj4gPtXy/mY1567wqlMYEhogDAWhJp7StJbO6kKG6Uj/ILfklbLNtG/dV8axjp8LsgdiqLlaKWF6q1YteGb9tFEssS2/n+vXUuJYslYkO4eXaYuhmI49t4pcEdOz6g9CBzieRAOUKSwzJFVbM6u6EKh1kXfkKMzUuEit6yYsTw9T7pPPot21HlCKv+Ri2qiQ0cJOpuhGiMar8EG9vk+tjiDhh1ooMkU9tTZItApT569C7/vepar3mCUDH9U2UqS4ZOgt3cpxma2YU3VS1EchcJLecSRg5vXSOMOxTp+mQ2HRoXjsIQlCMGEAqIjWnkql8CU9bTsks/P2wV+MJJ68Qh65j3zqeifD+oIYskfoWe+tDSNLn5BNXqTtD8WxNhE1H2KW+XQmHWMH4swBjMohhWvGRBDPN/IL7O6snzyfUqnHQmsF7dG8gJBCzYUG1pDj87PIq0kayiKdJXatuoPl8CjLgdGuYYiGRxLh7Qk6U31MP2EJh+n0Y8rcAj3m9WdqBbzfh3H/0JoC5TCof0nGO/VNMnUuca13ksP6vrJmMEw2XNZTy6uSWGh5lBxlLLok5ZDySeNbft+JnkOGxakkMm9Ec+/HGjpNApVEqepuJF/wgUW8AF+v7BDEPw0UglA45eA66D2Hnrgmz57hNepaNjzFumbptKm46tCU2NM6S3CRc51NwIJLisUH9V6QnR6ST/ea2wnqkFKH5F6PpZ8T0QxnScgZk6HXdmUKGhLRZnNaX6aE8rivLEU+b4NP2l6Q72cZc+vOJcWOVCnaPaVcIb+KKZFGMNlzhVb5dO9cn/bZJkPUMeU0iuDG9g1zO62RzY2l7qFUU2XHCn3kLTLakWfqziC6JxX3URmEzN3nhmOoyBSwC03KwIrvUGq67pDeLtGbkF6S3pOUTxn8XcoRDt8qHOEi0BjUZlSKNZ7/oeP3kdqcrHtw6Jm5CL6ETiSfdRMCR9ZNaOxw6JzQrgETT7wmSUqdrkY5qmWQTuv9yOoFCOdhS1WcJoaVY0DJzeo6Jj1Ip9WM1QQy9GraJ7nU8fmzMgyk7Fvtr1Wam0VBeZotlNMU20D6SJ6AXq9nPlIZ66Js2irIZYzjHCLy0nvmJPYeDFIcyMJ5XT4nOWpcMYhSpv4dyV0H4tDqFSCjou8p3ClouvPf7b51D4+NoiPpMq6p8AwvvB4e45RzRxYlR77G+Nz7KFyyKwXIGNjL2IEhYCKQHWehe1dntL4mO7nkjSyvm/IVke0aV3XKKgsac8hQCWfe95hztQRokD8RF8OGrBdQ6IozY2pZBZ8NrXCj7eYSn8uqx7TiQhxdT888Z9ZqbDt9kN5IN5rR0z0KfHt2bFcoFHuk0HLppsbcdLuvZqkLRKQj14V6lVfuzqjdQ/eZXo8E8KhXWoUGwurW5lG8IqWmxBiTlrXrHZ2AiuvKE0mD+qLz83PLhigpPQPyxKoV6IIN2pemBDnJ4BYsPSHyR16v8s8zN58Wi0AP4lfCI+7NQ2Rg+CgAdg0T15BlvGOp5/rCOKWWfUjFW5u2UL5mFOMs5eXmcGYTDHzWCuU4deCndAUDPKfTNofmWMVG3hS3GTUV8Pi2QzSxKcfuM5ZrX/NNg0X9cZOHo67kg6tayCO+xkoPwXi9agmCV4rjMG0tE6G0dWY2JmUifgc0jGnASxfTUXptsKrTqI1k7X/deWnDVehFHcmNqHmOHGe83ObRDHX+nU5OnBcqtGzPeDGzSG0T5SkDI4IYpnM94XIULQRPsUSNU17bc51zWJTFKsgY7e37RkTW9yfEZiYheA2DnkchpTNt7jRWMhwNTBHCidjaM8yaDscwDeJLYjwTNqUsUgLl2GcqV1b16SntTlJP8eH0vEZCby0y55+gIu/hu3sGo00ly1OwHEffIGnPiviMS7MS1Z0nNyV3Qz6PpNSB8qXxbmhjUinTrCm9KUPQORHUJklZGFL2GnsikITOlvYePrORi0rW+2bSOmShnA62uYzgwk0pGWqtK3RRmNq5knrimOZa9RbZiDmNX/fJO5OfxnEvw8Hru26UBjGyQSqfJk/SOLDMYjhXPcOVGk7IbWtGZjKlbQAOeR0Zs7j+qPvACw3JCW9dhqi15pGNRG276IBGzDXHQJQjK4+1B8vXVEoeGGLj1WgWXVm6QJxqa2EoPCfkLNpwjr0V+rTjwIJkyo1DYCiF7fnR7hnK6DiI19r1EgM1I9U5asvPwC1z+bXwVYhj7VvxedTi6j0KvGRWqMBszRhQiGwnQ5QMEy9lx6RmoIEMQUqGSAWOD1nKIq6mugYU/M778WdnqCyvmQ+lTtmjbbj2OY1u6hxC54pmm5U2b/lgeNXQVHBjRFtIRKEH++rZFugyLKnxpzg0EAeqgEwb34AsvOrhsu2uUdftDwmPP5qB5rM0mZYjTPS8k5mM29iJMDkvl+HhZ3WYMXW6RrUPQfr6AGreG/+LjEfIcIUKAPvBvK5/0uGs12gpWMhBwtiCQv0s1L8SgFl4OWfXn+QbtNQ+oUKaOPx1BKioJy1nWaMu/PK4vNp24HkGLsxQsdUB+exVnwgWcgC7RxKE51M3qvS+I2B4KkfGmLXpd6SZoUglLYQhSEuXTNrZBwDwQxF4ItDmKeA6Ds6H+qaxLAkmeUfG2n3mg4G6kYs6kmL+67vtkvKAWnR4HbvOtnZID5JoSxDaQBLrgIr/PY1ez9okuw7LdocBwTUuHdbzBr5USanp8zq7bAmrJG3Nc0cUer2vGgJ6X20jb5mY3kZPAvJmCE0GMX+sOZz2Gjpa2NKAqk9oHfbylBl6Vit1KI7Ab4eL5SCF7lQ1LeMOhZ0z5Vy1PjpTozRyGREnKZnk8GC1aQsPFc7MrXq61F7e4Ggp9fInaX6EdswRRVnqwRnhzIJskpGPLyxoHwOIuDWrCFOASE9bGRSgVik8WT0+LixZGpDOYXhMdLrDzrZi63+0xBJywnDmzRNSWirUvp7ASEgq1cT7D895do5m6Dj54Gdn9HxUvw8ZrMRxpdpNEVshk7yILXWwy2ig+qGk9KD6vZQbPvO5sT4rq0J9bt/nMJK4Qtu0WhcDWjYoy4cbbI/8vKcMAcD0bA03DFswPRoddQL7bPf2GMySWbCsONUK2sDcLsaBOKE6lPG25uCqfqMK4DLMS5KvkZBNpqo98ezZCkSxYCc9m8HsBlSZrjTqaV3QMYy+35HVnquIOiTXPPWwbfEPu7l3GQK2DJ5eJe+TTy3j3mQf1TJKqrWxlFvIUM8uoWO0ZnptYCjEqDw4oGKbIjfDoobnH1TmRqDgDDklf5NQvdqQVSEPsKu6zKyJFqVSr1L8/X1K8XIT6F7pHeMzYxylhc352p4g0sZN75JjLc80rA7p9p+qZ9D8OWpTXUONWzJswVMay/xMI5QtF5OnIc9+RvqZG0cQVgQb8j71q0KAkqvGrHtC/EIzBiWzbviQ84m1LplS+uVZwXBN90rAR4hfV4E8cX4+5RhE8+1lMOv7JiQqCN9I5lyrptu5jstueyusrYHyRas90jS0xqNre8mm7t+fgI68Ro29yrx7H4yuiyNDD45PxgMak2O3z4jYNaYx1jMybGh9J0NDg3pY1RIuG/UqL5v9C1RtyJr9rXXM9glzHaclnOpZu1lQU52O8rw+DJ2DCOi97Qe5g411zTr9p7/Ke1dYIPJUlZIheI0zQ5HhDULrGqxV2ByqdCsY7rwOyd1ti3z+dgos8jbh4boMM90n7qGXcqs2xNVclsvTPT8qbZeeTMtoBRcTIhOZlRdF85JnmPsmm/2R+fAwmUWi0uyu4TOpKyGTaNJTjxWoxdtKzG3zRb3GAToWzUlRrw6UvwhiyqhdO5BjZOXiJaGLcj4KJfJ5H/Ty0pORHhu5AXcpXK29QFkiPZ2tMLRu0sh4372u2dAIUg85FkP0kuFzUN0n95q6b9c6Cc3qZgo73VYS7epcJzJfvBeR0ObI57agHvlQelC6IUPvYJ2FNTa5Uof8cJI+VilNrrVOnvq27Ra40AFKMK2/QS5AcgeEwFSGIPVGjWFQqHNGepKLtXseQwKNtToiN1bd0+P2yjq0zTQTpejpacHfFFTsim8u7zmY4Wnk0CgOJ2oHlrxd3jM3I2XYqzql3OhKgoDrAJRyUwow5Q+PkKrByHz4uNR9zgwv84cWKsis0+jToIcETa+sT1Mca4YzU77SoREeu4x/33h7D5Ae0D30MIleoQYZ5mUnizBore2b5pxKPwFWNzbKKsPUyuSU/KuQzZpugkagCqkw2Us2EQ1/dJJ40zNEDtABQrT0N85UZ+oW2SbA44XQKRnsOlYBCDmGjg2L44TxXa6HHjSllLJaOUY+O/TaKaPcAxSUzkBx3DG3vSZNjQAAIABJREFUjcgCWy5YNEJVekgWodeSi+CaebEeQ/ailUwHmU6qHrjWcZ3Z8toZY8Fyg3aPmVGH1E49OMUBqBUcUJCL3nssa3pLo8CyTl/Kb+qNKK/B+aIdKBpI7wZMEmgzPU3pHlFCCr8jDBXFeN5PCu/0VMl5uDa20pzMj2sdyA3UFdptrMuw0soVHgDK2lRFqiB5510UhvCBUUCUhpOvkcG2NgbJh9JIZctNrI0Ppr2h5sHy0HWqWR7c1Vym8VRlUDlvlAHItn8z5uz8kOab+kSuQIVknTOR4YY2NolUQXeDMmNIFFlPK9MYZr2ea6geshU6ZYrSSxeRfyjTRFIohARVPCu7x4OZntJpRuCUzgRNji3Nr/MrKUPyj0TRa7fsMZI9eRZOu9JOcM+L98pK43dl/apird7D9Gh7qK7SaXCKhOT/U0ZZUp0Kvey/L2WfMhorEQgn3kg/oSQJcLoeO1dQMUecA494Otq9KQ5lXn0oPtTm5sBVnXoWhsoAoP07Qwf9eHk/n62X5yRI81JOfaZvvnwoLvI+xU0I+RByeIVgMe/y6kUMyquV185Es8cmBqyIaXl0oYREfGqTt+S8c32pmEVuz/a+vKKIOS1NH3OrApZMVZ9DolHtCjyvU6GVdKvXutRd0MZbCDAMQdNzn3kgz2fjwRRmaKzaQ7PQ4ExZawpbfTf3jzgHIRXkd9LIQDyM7T6X+pzFiXJAlEE6Xc977mSICNdGkWrMzxpz3WgkWP6OGjyA7HjVYHpu9GzsobMTfASeagcIu3yLcxX5b5078ajdn9sBdW5gw9xOCBkP9Xn+Ox60or6JM4ulwN9lYGrDohZPZK1ai51RlCKdRPjGQlx51zvhR77/q3H5JccJqbPegpskSc9umNNhbG0sJcoyvjybMSWHrUFmznE7hfvEox/9YPzjb30w1BQoZbOd5mfcZzzoKdeEMpqHei3lreuHDJdzx/iOJ34ZrjgH+C6sdHzR/e+Oxz7qvjn+pzz5anzL37t/GSovNHCWPAbD3X3NTxGjqhkI2909O9drbjB6gV3bABm0ObOnQ3XCUmMbzfVwRmdLzsEfUGaph6eRjkw5hX7PJsf+rFafp7y+MiezNqr0LEOfFjumzmH3ntGJVaEgUu+CSD9KfTVYZppM301iM2RYPWh1H9/JED4xJhVpHi6WYuXGq40cQgNUdBUdgny34NnVKa1zWbT9jQWdOOh+WInfqRx5vbb/46VobDoqRYQD/enm+VSx9p3u2aPRRwldRsU5R/gWRGbbePNwAp+neOLjH4r/6ckPxzd+5T35mp4Mddp+14bfUk5wJ/mkWJ1eUxuUdRaWMmjckYaZHaZCvne96grc5x6X7w1dbiBjXNzl2TxJkyHqCpCj8DlxfPll+KmnfwPuetmylyUMj7j6/njqUx6W8rvXva7EPa66A1TA5WcN+3bAPJyEM9i2kN3hBH6ITeib9C/+fsyjH4S73fEI1Z1KfSkYyjQjX3JuML8Z/dvrguRa37X+2al7oBV8dZ2c+XuXYT+6P4z9WrUeXt93dUHrhrW91+UHnymXST2UvOZGGW4HzMOF+F6TYTypD21NZvEsUgUhkNnCQMpmtZxU5f6n+goq/disXv27F5IQLilvrM/vikN0mGkQvslKLkEoNTUtT8y28oJWQ/dQnQTCGEAEa4s3cyUEWa2kkW/Ti3SSCm3xOR+FVrV5BjCAsR7jyY97MF76mg/gyY//MvzRn34YIknDgTQZchdVqbojSUXf9jLk3KrgSjHsPvUcBTnIcOjFL74GlbpUWBb9ExR/hpemVymCg/ML2RdydP6lCk15uJnfy8OG6IfDgF99zqtCR4bO06DWDITpI87IBNm4wE1xv/iuMNA2Vjzte74WP/ehj+CzN5xAZHhxZygZisi+nQyrZqJS+RA+KXkxPZ4EuvOchBpR24LRuozFdUaVWKOuX3OmEZJec+354ZAP389wuWVMupHz5oiDt9KzT7aSIccgRDKVmdLeIKqpsnSSwq4MovYQymAAvsZzKIvxTBIo903xCrXZRpFG0EZq5JMIGlngNFvdKOjfLYZXDOPcAFLKfps+EUN5AZGhjbRLPmOMbL6SSiOir8V6lYWgsmSBD5loKeCMlu8Pe8SDcPnpzfjV578ZL/rN78Hf+YJL8aFPnU+D8cyf/U68/mVvx7d+21fiK770Hrjphlvwn17wZrz3Y7fix37g0fiS+1+Jz193M37j+W/Cq/78b2NKY+B7/uFX4esf9T/gC666Az7/+Vvwwj94G176xg8BcDzt+x6Nr3nYvVIgDuCtb/oAnvcH78aTv/0r8cA7Op71/LfBYfiXP/MUvP7l1+DxT3wEHvWwe2E7PcWf/ZcP4t//5ptx4TSU/Mu+/L74oac+Clfd6Rx8AucvHjDnxO+/6O142Z/+dRmO/pstQFNKhaPpbQ34J//ksbj4sY/jP7/yg7Ax8Es//w/w27/1Rnzf9z4aD3nAXfH562/B7/7en+P/e/1fh0FYJp76j78W3/KYB+HOlx/js5+7Ga969V/iD/7kw/g3P/nNeNA9L8PP/otvw/mLG37vhX+OV731I7jjne+Ipz/t6/A1D78XttMDXveG9+HXf/canByAcXSEX/6578AvPOsV+F9+4LH4qofdE7/xvNfgha/+UKyjiOPUSS/9arq+49S0sdPYi4zkhoOcSzjSbqBqw3OPsFkPoBaQJFLFoUnhXbyS0pjiNsTFFAJwnMSG137iU89keLMKOpEWi7PszL5UaNTXG7DVsNSzYNAJJEAVZLLASXgli+tpLXepIHc+jEc7XBfsh5q8BLyzObR8E21DK7QJSGQuwjIs+OQhLsVjSrW5n8b3WXugWvkY5VnrSg+Z6dM9ZE0iLqAO4Bue8sSH4lWvex9uvvEWvPGaj+PJj3swnv0770wlvN99r8JP//Bj8W+f/Wr827+5Dn/vMQ/Fz/7YE/C3116PX/zV1+FDH70Rj//mR+Bn/rfH45p3/yauv+0AbBPnb70Nz/4Pr8ZHPnkTHvU1X4Jn/vg34y/f8xv4yPWneNGL34ZXvuIcAOCyO94Bv/xzT8EnPnEd4I4rr7oM974zlcAn7nOfK/GMH38cnvV/vR7P/uXX4O73vBK/8MxvxT/8+HX47T96H85dfin+z2c8Eb/y7D/Gq97yYdztC67Cc5/9XXjOv38ZXn/NJ1DwHZR9KPe54wWXnhNiCHR4vKp4J9Lv97jHnXH+ts+nIX7gA++JZ/zIY/F//Ic34EMfuwVXf8X98bM/8i245aaX4LVv/wge94Sr8a1f9YX4F//6xfjcjae43/2uwiV2wOmt5/Erv/5n+Ornfjee89zX4G8/dQE33XQey3KEn/9XT8HnP/xR/MCPvgDnLr8c//KnnogfHo5nPz8Q1gMfeHf83P/+LXjZy9+F5z7v9bj55ttKP7xxFk0nk5OV9/c4mJV+zM/E9qq6Bd/LbYc0oA4UmlAYOef+39ItF8kuRJEKy33SiEwXUhIhLcKSXzrT3czZV9UsLjmUhfRW0dl2SNaKMCO47kjKZE9VLMLfUbFSXKvXKtQpPO8bah8Eod7Rcy0iLip7phCnPpvKBwC2ROw/9F6VoJd30CLrbwqjF/DonD8teZpHZVvSKDFObIywmWeHqiuuvAu+/uovwNOe80fwOfHy174fP/+Dj8JzXvBOXDwg5/3a1/4F3vKXnwAceOXL34H/9fu+Fq951Tvx7g98Fu4TL/7Dd+DpT30k7nfPO+C6v7oBMOD3X/yOHPNrX/2X+GdP/Rrc/z53xEeuuw433nAeN954ETYW/MzTvgHvetN78Yo3fSRlYEBWmRuAN77+fXjdW64FYLj5Q5/Gq//Lh/GlX3x3mL0f9/2ie+LS09vw+rd+BHNzfOZTN+Ca934GX/qAu+I1b/t4KmyXoZnhuc/5/jOhGbAsCz70/g/Ts+nsA3ka2pGXvORteMd7PwkY8IbXvwcPe9h98ZRv/lK85q3X4orLz+HC+Yv4xKdvwvmLE+95z/lEp5/89E1wAJ/97E34xKfOA3B82dUPxIPvcYQn/9Sf4JYLG/C5W/G8F7wd/+7pj8Sv/s7bceoOt4G3//n78Xuv/ECtbwshwvDz+b25Xc4iX3Ee+r4yEns9hMSRWZDcc4hyFaEN7vtMeTPMNYWjdKC9WbEj7pFoZdYBQCBJWFPTYz51baAMeu/14iqTYIgHn20f7GG8K2x0YFUcnKlLzTG/NHKCuzr/9Dot1URCKbgmpvgUDijLkYfQJOQWG9moMJrnR2Y/H5GwrDpAl01R+kvQK+6t6r4YqxBHPyCl0KmZ7zQOo1l6Kgo1/wmPeyjm+Qt47OMfgcfCsBwd4bK7XoVHX31vbrT4+ehHr0ceoZ6Ok4sbPv6pG2gUDX56wOl0rGu1P3vIQ74Qj3rEfXHVnS+FmeGKS9lrMREV8A3f9HB85f0vw/f84EswNfc5K4RiUduHr72+jPIwXDh/AeudAwLfcN3NWO9wKe52p2N87LrzMAPufY/L8WfX3FJK616KxjX/oR/+bVx7/UnJEMDf/7ZH4nEPuyq9o36q/Bz48LXXFecE4H0f+DS+6TsfgGGGV73yL/CYr3wSfu/Xn4qXvup9+OPX/Fd88nO3wpExc/Pgji9+4D2wbYan/9Ovz3tdcZfLcdkd74A7XjrwuQshp2veeS0UVmQ9TdMpQfyE9EqR65xMykG8ViBZ1UlURbCXIYEhwoQFRYZOAgmGbdkHRgY5Jdb4kPrpGZEsBjTj2aqSsbKZuha/VM5TBqvxR2HQqqYkjZD4E0poBZUrfxgjqTQ2hLk2T1smM//bv98JUQ4ki3Ya0tD3s1w21XEfV/Vafq9bc9JOg3IaUFHVgu0glXgGJPcwywBsKsyiVW/Go4bpKVxZbcDw5Mc/GO9+7ydwlztdmovwvg9+Fk9+wkPwmrd+PD3HPBRqkdGZDIvC69bjGOHAP/rex+C7vvGL8Nv/79vxrnd/GIc58HVf9+BUeDhwt3tdhZ942iPxr575B7jxtkPGzYLKHWltp72JTHlLuOMzH/0Ufuflf4VffdZ34y3v+gjufZ+7Ybv+c/ijN/4tZTTrvm2db77lPG688aTet4HzFw7c2A6g+j/kGuifc0vPN7dJKOy4+YYb8c9/4gV4+MPvj29/0pfjPz/37+I//sdX44Wv/EBTTaUbJ44Ww623XMD7PvDJnVF/y59/EDedP8DGMQDg9CRSmKmLmfJtTiiRWKGz2ICM9WcYkP6O/EqA4YL60vFscpxeOz9Qa5FoN9Br7be6Thg41YQISUQRYtU5ESVTNp738YaOpX0RisR+NhgKzRQA4BwyQxMZunUX/4TEYFgwzJEVmzYwjY8U5JTluaxZ1UQnycCHhc1NZ9Zgmr7X5ehsiDNzYUQspcC9rifhy9LyG9CBGm/nKcryyvgAngfjClHpNkG5WEA2ehllIr7ky++P+14B/NAvvBI3XTjNasf7Peg++J1ffDK+8Ko/wceuP6GgqjuSnu+Q1n+0G5rBxhG+41sfiuf/2ivwkj/5MOCO5fgY61Gx62NZ8TM/8QS8+qVvx9ve/9md+pUYRcYhN1cci+8HwUImn7/hVlzz9r/Gq/70b3HDDe/CtR+/EZOIQZC3E3OQWplBDXwkV9PcEk3UoT8DcK973xn2gRv4/QUP+KKr8MlP3hQrRsT37ndfi3e/61o8+nEPxzP/6WPwklf/FXReZPB5MoDhI5+4EZfdYcHr3/DfcOEQlZV5aheGcVyeVnqcJ0k1PyIBT32yOijsE9WMmIbfVbpPBzQnspWCvoa6bvJbGE1/xX8Z+qHD+GjrGsbnghhD7blDayHTIWNmUVo+bKEfrUdCKpOTD+y2OAm82cBYjuJaEyiuriMLZUgHgAVDsUvUTlS9Q7GsVaUGZ6gx2+MGlftNKKwCKRX4VD+CLIBhMYtgdX8MXC/gqs/o+4f99/o91MiW4c7M69WDY+HORh5VD+LqTZGf9f14M+arGoG//4SH4A2vfw9uuhC1FLrnh//bR/Cea2/Bkx77oFZspZizE2NFru2OiM8Dbr7lBF947zvB5oZlAf7Rd38V7niO1t0d3/ldX4O7rxfwvBe+E0frwLoAq7U1pHLnk7PQal+E+DimuZ3iMV/7IFz/+VtxenqCyy47h/ve63IMzCpo64VJ8oS3k9Mh59Z/B5x6Ev/+H5/yd3G3Ox3B54b7fdEX4Dse98V45eveD/cN97vvlbjbnc+xwGpiHcCF2y5iumOeXMCNt2148APuFkbDDNe8+QP4/LwEP/r9j8RllxgME1dcfgke8sV3R+890gv60mhSb9XUpR6n2YuqJn9vNUBNh3R+Ym6nO12Ez3iNcpsqIPR6+LX2VD4lre3B0rPaf9prnUjNIkftmfa9Pm7pZiFTtWK0tnfaWnd7ALBO4wDHjDBkZLkwII5iYsTrfE1HYGV6DbKEW7OgSI8Uzyzm06EhiMXmNsO56BNjnIuB6utjCStolc6UzR627mIyt3htqh7eFKtX3JiH82IQlf1oee6ynizLpSM1W4I1hwO2YIwVx5dehoc+4C74xX/3xujbYHPnSV780r/AP3j0fbH8/ntx8eIptkmvS/FevHjAnBaPRAAAW3DhwincQ96/9rw/wzN//LH4xid8BWCGV7/inXjtWz8Gx4IxjvDtT3oorjqe+N3/+2mJpN7zzr/GM571Rmyb4/TUsYxjAIaTkwO2OfhU8BDw4eA4OTiGLTh32R3wyU9cj2950tX4uq9/CGwMXHXl5fjY33wSP/KMl+LmCxscW/Tq8PjOhQsh63jawYRS1ds2cfFkYuHZg9PTDYfDjDXjIvzJm6/Fr/3K92IdhisuO8bLXvpW/OEbrsXAwAO/5L74yR/4Kpy/7SImDH56gp//pddissPZb/0/b8c//9En4Xu+7zxe9MI34Xdf8UH85DP+ED/9Y4/FH73galw42XDJuQWve9W78P4PfAZGuYId4EKX2IHLPPSFLL8eJA2FBknmLojHfqxQjK/6EOnR0KG82BBwdz7fg4jXdeaKYYw1hcyeICN10LK2CfvwRIhlOtFBO0RnGnaEF2brbl+aexGVEGdU1Z4VJimZUOdBktvZBuzLHvnj5229yyX8dG7QHgroidtDXau9NlRtTA2GILcf/MnikQaPYZjzJE44kgsx2L6IB0ihy7vvCsFkkNqjCvLkqiCamPw2tyQ5z4QmvRDHfaOSFJIx9sUo8tcQDVM0ZhqNbHy7ny8gDoahXSIXRxVeGY6OF1x5pzvg5ptvxW3nTzEW5uSzGU+FE3kMHkB/xOLQU9Ktjm4r3675//TPPAWnn/w4fum338GxGI4vOYfnP+9/xn96zsvwyrd8fCfrjGuVzXKRgZ6K2eUbMjyCLQv+8EU/iH/zE7+Fd/zNzbjqystw6y0XcOv503AsPKNzdDRwlztfhu1wwA03XsTG6lltsMsuuwSXXXqM666/GdNVuLThjldcikvODdx8ywluO39yZowKZZXFUDezNWXfdaGK5oCxHOdDeWotdQhxrWP4/cfnzill7U7O4/Y/mYnJSCXOOMnDjzxXo+u1cF564LUmYyyYc+P30OZJA2Zr7r3QwzoW34++d731ww0X197nsQ6zzCQ4k6AiPOkXVaRfAkFZTgcyMTknbIh8kXXjZwSTQGnlJhslDI4pn7+ZcNLycNVQkVjbpDqNZxRyhY1KW/E6rQt2CmpOHs1WWIY8oAYRpBlVaNNPXbZeb2cZQE6mvMrMRU/Y5xtOL058+jM38HVgY7n4GBVjl1Gb6blrjRv8N6AawYpUCwj8oPvfHS96wzXw1k19jIGjI8Mtt54ktEWmtKsCILkjq3nuGufGZFCkcPz7cHqCz3xmS8MiZXafuHjhFJ/+zIFevQx4oDzDrbecx623XMh7KON140234UZIARFduqSnua6sTsx14hhab5A69GeU0WFnYLSjo1/m2I0t0HcIZJcRcmWoHNYzh5DIaWTVBlFKqk77Cvcg8hjkkXiqViESVJK+QUmHOFRI8l6OygE92CnWTXKznHfKPbmnGPMa3lceuDaoz1MKfYFPD0tka/aFUHjQU091E0AFXeJgfQbBBJNHiHtgFDfgcBghb0B0KwOj8l/z+F4uNA/26PSkIJy1GNWqlbqUtq6d+4uvR9gx5ykWG5h+4IJsMeyMJQOO58lVKUczOs4H2ozlqBaVaAhYarHOjsnbWOGAc+5oHkpdqOdpIA4ZSmYixlhj/Xru3hZMEWHzFH/48nfjnz39m/CFf+e/4robz+PKK6/AY77uQfjgO96PN//lJ/iAGRp7hU3yNJnjbik3ebEB+DxgzgOWxTAnjYwOchlVninIbCQko8s1kz65n8bnqPBznkbXskF5aBF3Muwe3+HsrxHNjiYJ/FivuZ2mQVf6OWR4FOsrzgxEZ/MABzc4VQdtX+goerzJMu7eG3MnO+qnKiylR5Sh+xZl8Y0zCgslAydDPZHH3/N1GRfVVLDDlkW7wjGOmgwZbjciNZeUBnK5+72/+hljvXxV/FLxLTeuial2stH96UwauNp2WXohWbJdnws0Kwx9ptrgAWDdvdj2sGpCGXr8oay3WPWULrQRveKthJW+v55rgdHu5VCHaR13r6SYRTszng2I60R2aIwjVOuyBWO07MXYt4AbOtXbISnjTfFAyJqPFt4lt4KSc2hL9U+AMjZo/T7Otg8snuED7/8o3voXn8Bd7nwHXHaHI9xw/U140Yvehhf+8fsxcy8JlrbYPF/XelqumeZYOhQy3LYN733vR3HrRd/pmbW/hymOXpoeWr6GlvVSW7iUE8OslIFk2D+TY6twUD8VHpa+qWBpL0OmMZW65736eY5+ulM6XmUAZyF+rSsX7vYybKEl8p4LdUt7IBoEGyzbSKYMuTbaWxqnskuF5PXx/V6CDWBe3OwhX/HD52298hJ5n0hTIhqlMq4b46geqGpA5p+FMOQtW1yVzWUo7OQJ2ibJhwonF6Fa+0a55MLUWXxXmGSGMc5F5sMsFUX8h1BBCJ2HhBJ2hWQcnkSuGgk7syQ2jui5R208Qs3dA5FRhklCdjjmdpJeplLBVCbFim2OcTJRct2w/7FM0Uq502MkZ+ElR7ZC1AOYAWTuP0lgop2xHEPcRG00ypmczV5xS+HNRqQUc1099WPOQ1w7ZViKCCsZ6nscJJ3CyvkdSi9zXqdhLHq7R3Fb8rKSYa7L2I/f6gxRpYeRSDg+sjQdrbMw4rMmuTJXkZaN/Hx3cDG+QgC1jsGt9HUX6tC9A3Wthcq1DjDKasJkzIX9bAn0NY5Chj0TZ0Gkb0QWxT0BRaiOXA6N2w+fv8gjdhUvqwArjDEnpE0AKpG3RW78xSS5UqRXPRJPitVRhScy8Ob5dR+TTu0EFFyEGOrZrlvopFDDaHPQbQsCAsgH/PTTnqksOd/Ktcf5kub1HRChGjLU7yQG0/DR6NHzw+NhxAKKmeFJEqptSq2zpJCMeRmngMmHvLeUKWUgKoHKkAcEu7yTrCsOJK5T52dqJKjPKPwo2MGriutQj9Eo9NLJzrwWIXDOaU74aOm+DPOd92rrLESZnc3YET7DPd1mpLyUCUgHMIXOvDmBLeWyRwTW7qsaCdZyOMoZJsIG50Xdt3YpoOo6oPC1EKOQR7wbnFA+DIgoQWFMfKU3KiqdLTmO9l2hh169PQgGZEQbEWwDK9zryUOw2jxg0Ucqu/4bRkAbsl6PzxsVLAtpbA279//39abNtm7XWdgz37XOVWtJ5iJbliwDDkkFynRxugpVcdxUqFAUf4OflL+RokI+pKtKydhQAgwCTAWbCCRjI1m6lu6VJd179pqDD2M8zVznOPvaOnuv9b6zGXP03ZRzZRa4X1rt5Nj8XRpGRiwmmoIuHruteQ6tlG4iAJNvyGGzDqViD6MhuOWfkfqItQYDQ3EPthtl9g4CJQwBEr21CiI80CbNrtegNoRhEhez5gTzYIJYYp40lbB4R2bhmjChnchsWOR9z+y4LfoArNqTkKWpKPOvDrhyBSJwEeycw7rkQwpFf/Z+xc13ABPViNQiUMGTs/k3MtRrLWzykmWBci3DUOukmZDwY6craRkMzzPhcMGZm33G1+2OXdWfCobwGW2ar5dxrClwiDvOEks+wIVLdUcAr1PwKip25D4Z3dRnJb6HSf8GE+es1ULSeG/4gg5z0eb4ibAm3VtScCFvUnZIJRx8lZoFvbgBeFitaW1jvNY7i8/WvPvQBTsMwTbiFnQ1IuO9oQ7TCw2UmsmyVLpmXIbVajSkvm6+JdrW7de0a53yLS/8EU6ixlB+h1GU3RcULZR6EqjFOb39ygRk4dv0GGBLOMJwwo2Ho2zOp8nsJpMFRen/0Jo6NVlY0d9NK33QXzHv53V1wCPGfaAkwQB7x0/4bJowclDeRnEprLlarxPejLBM9YZ8MhUSMBhUz2D8wXj4Udjj6Fv1wJ7u64Vxnk9W7GE6RDZjoaYp0tIZpVOvTcJIlFvc/y2IfyIP7Bs6PxQUvacNm3AlQXI0Hx7Wy5SE1JKr9tT7lByjZGrukWnNpWFtpls0v6ODPKNmBaCqu6Z1V3/SHl0LrXXzLtQapz9QuLfD7d7JU1JN7n04UmMnn2CNjbPtlNnSusYmlWQZWxO0pxAMabz79ZiuR9PHEQUc+RiTqQkyjpc5MFfsLdyh6xTXcM1xxvX9k5Da6KYxr4IpzG1dGEWWlxZXzX7HRLqu/pvD4WXs5gX6NHCdiTfXOCJ16c6oeHTWaR8XZcY43ygFBTPSlyUBGHrMGh55zNdBhLTrz/6lzk4Fmx3vPclDo9nhBSqhpllHqbacJLcLh1l68VKgBaz4vQbOlFq7hlD2pf1ISxo7/nZNQ+BZO6MmTExiZMzaBzWqa9ZMql/qadIwtTa094taIyTjIoOz+s91vLwBw/ZNMR9iT/f3bpOAdalr/nnipa5xAAAgAElEQVRPSDvHr2vyOQDQL3HJv7aUt0PnKuHRODs+kjFzZYrsB671amB8D1OjhSPzg651H38kk7MGNnSaUqOshft+ecH1atJHR23mPQRrXVMJOqmhNdlpe6MWw6ojCZmTMAgzjoU5mAag4/CPUTnD056K1mJFHkGKUZnY4Wg0k0T4p8atR10K1qyZsWzMdQGDgHtMmXp0r1m2MQuTo3sgeOyG1xYCK7RbAJvTspkt5F+Zw+RNXST0zF8ZtV+Vnop6pNStgbFh19qIn1/XDfVgM5+B2Ggk6RwjwRB2a1TnJc2C8+X6IFPjmlCkS4CmRH2/Pp6XFrF8xnu/btgqz+dqHaoKj0V7ewa+WLU8YUi0xFPiWfX1ghgThxpDK+mjWsufNOuZ9dKMJK7ot3WhSNxU19dqIUQncBnHOmpAfrQ1ki5dHu0Sc7ZFnMGUJvSCet3X2Wu1d0R8BwrUnl78ufwXG7teLCxgR2nvq+F2VWFfNTAMv8xYFhhRTwF9v26TOnrZZ8CIiDjhWu0hlV9hzm/Cc+TsDMtRpVZ7MYWjxgm1blh4jIlyw1pOorJj7y6A9pRLEngsRnFYVKtqa9lOPLMyr/aPTCiJ3uwlYFy6ZEbFUdfSYWRqrBDjos15jV9mH3tdq8BO2x1i3QO3cYaBduyttzV2c0uKiyuzJCQj550O1x1rb2xMlKrQjkvQY8FQGsvbB1bUYmg7L5iA1hVrDTONZ1wuDKMJ0iE8MgBGrFZLpkVHYiQFcU9gWPkeFcODpAt+NiQpqJVd9AVNScKsiWs4kH8tqDP2scZxUM7znfXYSWlU2RuGN7SjHjqDa84N9AksN5RZb8DQAs9RtVgvAKae05yuRb8BDBs52In3dLCSJVUXCjKyFntuMI5GJ5qGonJsE0g2pJyX5bGvdcd9P16w8Ho2PU7IoiYwhEkJfE0y0XDJPYU49uRTjRwtgjbASDx74BmKW8HFqDYuc9h1A+q1VCICgj+L7880hgzXX0/PZIXh+DeoBVHSjj3dUh8jnbro6Lq9EoKh9jigCpv2r0wCJlbNPvfrWONIJZpTu/8VYwy/j8PR3oM+35NEIy2r135752OolxfD67qpxBpU8tbCZ/78f4L3/83vNvMhLmuekbRV6HJynPPfPo7PfvlP4/tf/z3vg+ptebwO3S5pB489lwST8Vah7eeWmgP5WYxbzfXfnH/gdUFntmB/EJPTBEM54yFGyqJCzSfxyQzj08ktCRl+Af9OH9v19N0aWspubPT/kCkObMacVG2S5twBw07aavOeDCpxDQAesYatZC5on03j8rfsBbYLMG5luUdq/NUl6teYHvJEL2DHjU2LQBERkuhHZdLFJtJFoczQDOXRaVOsvOsMR19bt4fwRgVa01dj0cE1kmEyIxu4l+3W4bZ2BhGIEBJT3a/KSAXVzAELPcxFW7cg/w2BXhi4OUbPyAQZColsBYMjI1bEgg6w8WnwdxY5AU7q6ekf5OOGYRU++eU/i3f/8z+Hjz74Ae6f+gl8/19+DR/8/rda1dw9dkWuwWd+/s/ge//vb/ffGmvjY5/7Cbz84H3ULtzf/QJ+6i/8LP79V76Kj33uc/jwe38EAPj4F76I+zsvIkpGDUiAHI97UwSDESsSVNX4NFxuYPgvSWKIyOnLIt49DhgqXF1DOMKzB6iTtr9hC4ZNV6/B5kjtO6fdT9wmTqJV/iFEVX1SgIxjsAslyTFf5q4S1kpRUDY89t6tWQ+NkQk1HGJvtUJOmgGiaqI/A/MQuDI3gc7kHVh1nsdjrkfYeBaomn+H2aN+Fk1FzQToTJGKk/baaBmbxLMm3EPT5T6LHQBGEtFFZ+AACteF/VjzuQ/uWrzhajSMyxl3TqXl31MsM8eo4h2sTkCaVGhQcoXqycOsYoEcGTrXGEgdB3kmjT2pmfM8k7X8PfsOhDlELYeaBqCx2y4H3LRmeOG6jzNy5l4YpnfHT//iX8K/+1/+13j+httcZkzzhO3o1/UO1uz7ut9R04Rm7xe8+1f+Mr7967/ZCtF738V/+I0/xHW9wrt/+a/gD77yFSwsfPrLX8IP/vlXHWa84Nb1oWkystVwDQc6qA1JYYBZ9TybMAUZDmFy4Vo8MzJUBAyJz4CS4iKiQDwWYV7Eibulqt65BpdeZp67hGNvObKTL+ZuMPOXuUQXCuOQxTjza5IBr4ULtzY/yXQJo0UYDnxq0hYCJoPwQ3fDnCNaYg2OeMaI0DW+M6aiL/nkjENOo6h1w52SXioKG4lStRtgdDYdpWIBcp6QKMJWlGbBEFTn85+Vngu1P0IBk4E5i74NEhDYNG1WVEzuF/lKa71oXl8vUNMzI/Ljt/0aDtP2WvZRILdm/bNXOabMsHRAqEkgstPMBUOUrBFio/Py8ZGR9+mn11IjtSyBWt17rTUqpL1fJnDSjir7aAqf/ou/AHzv9/H+v/82AOALv/Y/4Pf/z/8Lrz7/RTw+/BG++Cu/hNqF23rB7/3fv47P/aW/hs/9Zz8PPF7wR//8n+Gzf/W/xHd/49fxp37xv8Fn/vzPYb/81/juP/4qPvapd/DdD34M3O74wi/999ivf4xP/NTn8c2/+/fw8joqPAO3qAkahtasJARk6hQWC+3orNRPP7/3R0O46eRuRDc+zPuTjTuIMM9bPW8YOsmPGgtrQ64qR/fmbHxGDofLJIgb1FC7W+kd2bDUDNeE3m0CcQ/Ko9G4zrwVG91kCuLUgkXVlubrs6DArFgnI2RmzhTEBHuha6Xuhe37F3gcVN1CQqosVw6ny3YQcG5iNswQIrefjjQ6czqMOE493WmxkFmRrn3wuMNMm4tPJaccjXM7+4lk1CQcUbBQK6vNeAwfSG88Cb/8bkU0J23RCYm6NDqZUF4UHAVe1imf4BWMtRKJADAdbRjgd//Fv8Gf+Zt/A9/6jX+AD7/3Ada64dNf/Gl853f/VTP864b7Ox0y/vSXv4yPfeaT+Prf/d+BAn7ub/9tXNeFD/7tN/Cpz76Db/39fwSshY998uPYL4Uf/N4f4Prxd/Ctf/avtOeqwk//9b+OP/qtr+JH772PL/zqr+H26sLLR2UzkR51mq9gZIJnwXTs0rkwi7Pp/ET+HjIa7Rww3MIr66k1OBgOccJVzsaFzGikZtBruU3H94VV7Bp3k2Oevq6F0fpadxceXtRypCtdE0KnxjW0JB+H9yAWWRTOaK2ELgP6FsBGNmNHx1iFh95N+FOINX2xGc5leAnX57zGvL6znT4/oDpD3k+ggcQxAFFqqyTC0v9zA1S/neY9o3L9817fKLYEWDsy6UwkAETdYEuxRp4VRFlS12qkvz3H1wlQxdzHK87EnmImI8NmzUT8c2HxMumJ6ZdWT1OHzMhwoT0p30qo5q0y3iYjL9PAXYSUmk3CcGHhg3/92/jR730DP/Mrv4wPfvuf4vtf/wPcX93w8lEjwu0n3sXjgz8CauGTX/w8/sP/839A950+Oi/gk1/6WfzxN7/Z897eAR5ty3/qZ7+IP/7dr2HVwu3Tfwr1w/exrnfw2Z//OeDDH+Nzn/g4Xt77Fl7/kCnSYxNPRmmfyew38jakXai3BL9ideSCurGL2d6BTArUO4x23LsVHQKuPJM5n16HlUPMtzRDxWoC73I8w9+mepWvpnAp+RBdOwGVh2PzfhlGk0CWwkOeh/VqGCNpYEm+rBGMChwI130Naac1GN/XNPNRgZoAT5M/cK5o/l24ty3mMnN7Q9vpuEb93fv19AOk/d2cVQUr25JBkmSX4uAuGIO8/t1w5aOJt88N64uOvWQAoRoN06lhFhcW6CglU2oGRdWr/RXt34DWSSYiD/AcOAHm8mlKvQdWpenQnnxqAxlHTxgy/VmqH1ZUpdLZ2306Vk2bN8GQxMLchmjCstxgpjuoPfDRB+/hG3/vf8Of/Vu/iu9/8w+xP/oBWIz0uf/0z+EH3/g69v4Ir94Bfvje93sX68J1K7y8fIRP/vRP4ru/8TXU3njn3c/jw2934+FP/OSn8N53vte/f+mL+ONvfB3r0z+BH33zd/Cd3/onePnRD2UnN5LZgb0EL+ZJTF1ItbnbWZg4zpqIm55+mo/rUdj1Glc62YHuAo+FtSbZb50l3YVsJMPMU6+LGak75mMeB9/h53s/Ju/D2bPAbebsuakVSkMfx/Se4j6FSQdG9r1kVfc4pw8Ny743cTtqnUr0Y3rAK43rcDGaLh8fjhYVNHD4ZV6jzEZQ9cCdkygWLZer04Q7nk0AXloYMBmPmMKu6bbEnPP8fjWkQXOEZos5rZlw6DTzYajez5Ebjx7rugV/RuxpSX1kFqU+40jirox1t6rawZQ1uRqBBKqK5Do4HrDwSmO6dRvAKMwut1rH4tqY+UopQelmp5/XO/NdfafKwsLHf+oLeP2993CnJgHg9qnP4Gf+u1/E7/zP/xDr/gl88gvvyrR597/6b/H+v/waFhZefeIdPD5srfDTX/5Z/PH/97XZM6XohU9/6afwna/8CxQ+gfunPov9oYUBGSfV7I0thzVVXrVqXET8qagU7GgeGFaY9+VkZwZxRqOINxFu1tkbsYRxDHnaVT1ynM/XmHiJX2XG1rkX4cSO87fGlGZ4n3Pv/9KQ1r5MN6Kz8d3Y5OG4S89n1itHvNatV0ZYC45Lv1/XO+gcnxs2XLnc57fQBaUBt1q4D7sDPcX6cr909ma1GtONQ+5xT6OTZpq5sTWewzit8Y9JQu662I9yiZjXhEPWmvqHSGhxyHIBqgRk4VP6JKDCmaWD3YcNxx+ZK3ssw0WUMffuEJjDsi3lmKtQgyjb6EYNZC1JFqcil+ZkhyPqDQzxtabO0nsyR4eiQVycv63+Fn7mV38VF6X56x/jW1/5TWC9g1ef/6v44i+/i/3hD/Gd3/wHePkIePXuT+Lbf/+r+PLf+B+xHxs//oNv4L3f+SYA4EffeR9f+rVfxnu/9Vu43TZ+9N0PgNr46Acf4ku/8kv4w3/4m9g/fB8vH74A+ADf+7ffxpf/p1/Dy4cf4ge/86/x/r/jxUR4guH0WK2yH23CjLiefUEjrR8MfzOsyu/GV9a64JgDND/3NEd6CRhGuLLYggDzu2GIpYwJEeO1LuwV4fXVCUwd7gRcNTxnIiHZyLyqDjqQ8IP3XCis3SZWDb53VHL8g+PAdpJUjfmyJiT7CHOIMKTztcQs1X4BI3znTDqStb3uqoYhBVnFmn7hF/7Oj67rcx83h24gd7447fyuy7jmLgbHuxHZco3NhxkSnOxQobFijqwuLdj+XwEc+HcsIdBzc9Sey15ttVKTFKNN+WYU4qg9GBPCTV3t8O0+Bo9QB7nvRGzme7zIRjTc7ExzZMU+Gsrw0l8VY07OSiSpuYVcxbtWL1sVtdc+4UEYKt+E/Fnh5op12xa3XV/n3M/ON8GwAobsT1ljwk4z3EH3c7+9Pof0ec5kuoZ5SvBT4nOvl/6WBnPA8MzL6f3cptvXO10/Akydz8vgwWu4VAHG3XXF+m0WuM8qBG+fi80Q4hSqYdT440CDzkgCyXsz/MNcwRSsLV4VQHp+BTldB/YM6bb563H3/v6HbbhVIBm5PMNdlLo1G5dWHLHwitwCCwmkHcoQV4lT0fkDc1tob2DKeCiUkyH5SsxDJEWvMp2o9CD3S217SQKtkziFIMH1xaBgH4f2zajPEmKumYew6B+HXbPsn+E8OW6XvfROswWCbEBi6/yVbeYpr7b7TRRVNEofXQw1RF4vWOuVFC6agXTGmdgS0VlbUYIBJEUNQ0fH5t9q/FFonj+KYKQpiRNGgNdBvBzTgDeKSYMkDq1heOIVs4ZJaJIfqB5RIpJO8WDgxAoxERm1s5+GMT2lUuPpu1KUgj6obRMnGVjgXIWEl9Bbxm/tB4NP6SQm/op++2xUF8PxB247/CStTSzxAQjvuKUec+I9PdglydvSaq1XsUBqGUZeHRhXl4eBAlNu2ZKPDMZSrVNOD6RcrZUUKDEfcMp5x4ZZJQfUWBolc4kE09wwCmwojVigVnRoUspY6ihzExeQdp9CcBgNYRnvJ5S5ppagufUDXam6PC/aJFtwGGsh1NdhqOlQk4akWpxyzouYcThX98sUeJ0+gRqk3fsxvSV5lpcQmfkr9iP1We2oTTBRxPlmQpwk5cCQuCfVv+e7qk1MdoEiE76mCxbzRm7rlSU2JgwZvx8EUkFUtcd2XwPTTIe2adhERCc1JfjGdQHZJxRY2Op9yvwewikZC6DogxhnMxCF3FP7Fn5SE7CmSiECOeI7/0a+PvmvEl8Gx9YNPND2HZpanU3L8KkOSczB+Nj/3lccEsQAzEAOdkCPquyzk9NZCp2miN7RTBwzUoWJAKrCnFL32RjkuLyUcSlHZeUVfTZXKDGpOkp9HruMz8uuRBH9kK4vtRs7wrn+7OieVdBdKZL4yfmHaJgBS7g2FI08VMoRTKPXeQv4Xzp4JjwpQxGNrHJ2zRpYgn/xDpfqMHHf1eI1Id5pSTdmGjWP0Ro4j8xYAKpElkZDxOdaR8tZtomtJ4a2ioXOqbFpBikSE94WbvLLYLxrTcWncwVQ4TzV/ohju2E6AoRFfp03cRmX5jzYM9QSe53jigDhOeiHCucnYs/6lTDk+dN/UBw9BFqUD1BQ2iwlDsdMIwzUwZ+nTEa7Yi18tqpDp3suKyaXwcJ0UH7VQcoByBUJOQY0ESUONEGkBdiOcnixYrwhFmnz29x/hSaAMDFQfXN07SDY/P8hXnQegVQ5Y9cgZeRfRIJWZ0gysSWamRBZmeux4mCDUN231NJf/UEq1xFOuOMnTJAC2LeCSC/GB8LAWhtD2zW3cW+U7xIZpLJl8DByKPeEkCLC7vg9z5YrTSKFYMgztCqPOZO5g5P+DZ3ojLeeTEfCbPwujLcQDt7Ts1lJQttIHw7zE6yZOc1bV0jIsW08qKsds3sRR0ew1FK3LsOHTu1e+2EGp/CgKQOHzNW9vWqO5KF1NsN+dPZnQM4zT/sARaj4LYXd9BFdrwSXFQzbJvW5nzvDJ5IKM+g1UuMSF7ZX2JzdUsIcuv/b2M77rzq/VZKXi9gaqJHgNGNfRJz5hj00KrSWlY5FIkh502zRFoXfBuIcxiFhEC3hFjk2d3bp7b58KTWOlFhAh96u2JM1noU1MX3L1POHyB4HVowsjSY2anY7pEZ1ZugXaxrZXNIAWNJNxlbS2wb5YOkoGCU8h+mLEce6XETXvUU3tbF5xGfTjLnXsHiqHi4kdIOA6jzGJeHbN9bMI9yisxDBMHTOZBpmvBSQcjKOfyCTEC/uZ10Tg7tUE7PL+H/mmZARXMD4oMgTDMPZ0MB4DeNwK8s+kzWLZxJkwlFukkM4bpCmK85pYRgScSc0vIXlJLPKkD1h2P/el7SNHcQbUq5oKw65DgJfWLCThz0MaVeVmAuzEdda00OBm+1jV+evIKLFsRHql2LQM99oCtckw/RztPW4/jMkSomstOBFNhAHAGtMq7wORkOsPc16tJf+l30sFdGJ3XnuEsw0HpmSDsuIcE3jYyKSQ3ZNlm+YeCSGeqhzGFcpRBltDWLM875g2Aim/BAxLiMPka+/oRTLLMUrYDuo+8wQOBol9GhrV8KQRDZUd8HwOWFIU4PMxo49V1Y38yQs7Q21QCOduL+o8dn7tiAVPq9rCG4JLgyjrymyTHPtfI/nVIIcM5F03oIR907zTk4AnbOiKHT8ji9P9Exa0qky7+RCZw1TQzUF3c0U+EX8LdXGXmo1xiFiI1RipHp9wH02SuKyqo9F6W7k0bjLKtvKQhw5sSaeTO+4NU8v4HAiEcjc3obd4sFMyoTFMcy0IOIkN6aZJqYQ47x1HbOAlTAUtBNoXAeO99I/pI5a4VehOn6GPOckI9rS5wDoEmehW4QthQuWgmQwDLXlj5jDk6lqOKzYA2Fg5nYwpWIUicso99CsfN9rsDTF8Uxvl+dNH1sJVmR2BbYe6LW0XT9mDBlT7SniirPbE2EpRj+0IP9CvHqCmQsged7O57HTc85gtLgejhqUQ+qOfgUTlcmK8acRzwgfuxf68WgtSMaJVfeONrCmPe3zh7gwsCZOe8eJP+mASYQgMTN5iiE/96XguywMcppzhhY51wOYC2a76Uv4DnRb+R4mGtWprHwVZ+29ZtbbYiFNvMf9Y+xTSwSghhjoQe+0dft8+lgeYmTWORx9MZhcSOUPDwwzkgQD0P2fQwBk6LKt+T0KrFx1AVFLU9v2BTxdb0AJ5PNNAZBMYwXCEhsBak9dsbnMoKrc6zX8Ud3kBYY/CioSI6KHIuL95Y3t58+zZpdJhL2/l/iuxByAjgi1zY+B+ZznJCPK97bj/NblhkT8fmgJevbZhCNBEx+DkQhGXTmdcFbS2dP59PKdd0La0Dp4vlMm4HMVRxAjP+kZKOzOxe5zdBy4KBVXQSodJZuxBhgC2lPb0J/vA5A1h7KuKIIalZDZZ0eS1XoFRx+uiWJck1WWTrY6mEBikyIxRMg6N07ioRRdgxQAkYPVgHvWQGQhV376EbMJGAbBNZH02LppinvZfjebvZiJGIbUCEqaFhkStObTD0IHIlVKE8aZSOXqxZ7GPU1MXL0mFoI1FNIpy7FLjJfMDMwrKHhdJ/UrOpUm5DGH5qVw4iJyTr9LOBlHXs8eyFr5VencHJWqeWeZYSVzrSZY4lbWLTkhjATczIP/YqXW6p4mNsGSRpg/VN5rEvIUAmrtivDxvODfY+2JW62J7iH3JxgM/LmWu7gXGGacjLpUuwg8mgCSLunFfoGdf5T8WamJWdw1SNPqD1Ug+zoA9+lcuNRQB9iqQTC6NjyWG+2kpBHhoO96CBU9pY5BTA48MLlsXlgbmbfkMW54dJRh7GK2MxtpZCQgDE9kUFJTOeT4bKIM9Oas07HMuoLwETFiEi3sMfAu0EdBibT0nZxnNCGo8BDSlKCxZmoMEGzYV4NMiRKdxGP3pBnRnEO9wLkwd50bYC2h4n+XxqMKnWeJZtzbiX1KcuJ3hKEcz8y8XMbnRdiYoDsHidWvrGJtwlsZLn+b1lP5NRn2DSn5UdsaIqgd8uXBIR5r5d5Jy/QxUTu0FkH8IOPkTe1YhLV/1jBbdszqTllsGPp0mJI0RduHrbkwwGN8wSqpbHttnFqIkaI3PBtlVSXHTscDG6DIwXOGnpKL5zV3ljqHO1KIJbQL+8+ZeCxOgg7mKGYiZx74NBNyIZXSkznTbJ/IevoRLMtBCcL1lUNuJ6YZ3pBJdfnz8P0IMw/JQim5NYZgmGe/AHdt4jBiB57zDSaAYEZcgnNvMq+nyDQ0nu/ShWCR+/E5Nt+64lOPmns1DjzDgn9GyDQ02mMMEZwWEIScZsBoepGvQnxRxCXqfXT25fd9tksww2ilLUBbW1zT4zZTEOjv6M5bFfMEHi1CaQPbTYHkCzokBGm2V9q3qMNt74+qOzmDMEAciTlj6njm3Wv58MiFTQhGiirMbVK+Is6x3nHWcM5AMgOwaYLjlw44JKt4lWspci7wkyLy3wE80DcCD5AkYalRkfFNYd0wM/lN9ON4NZu5EOSuzkT8G2taDr9ZA0pxxDEB+8wTho0wkN8ntJRDBSYROrLAOZLxNW2E5AWl07PU9Hzts+GyU31PhzJa+NSkzM+zeWMXBoZmq/ztFnt7WgVxobbMDK2Po1RJOea+jn8HtsS/dspnYtnbYOgzWrCGwbtXKAAOGilWaQO8m0SCiWbcvDcnPJ3UOvnuWatogn8I9xzGDSFZDpc3PWd05YRhDQyBRvU7tQTohcsTzuFck0lpDnFKxP6VUjTUu9LM4vJSj3iIMhUWIN/FBlvTaR0FEQ8Bf3ZGqhjD6v7ZBHWYGAEdx8v3me5v5gLQLHBkAg6bhaQ0E2VWnUCIdRDJMIU4IHO3hK50IL14+ET0McPAI+GJQLTlBe+QouWxemTnzZAoeE5pGvW6MhMx94i5jk+bCliPVpG5BVOBi7zSj4QuhiuUgzJ5qb2tLC6Ls5XO4pUYBsbN8x4WQ7pGe2BdSy37ElSUNzC7jsLFiNww27UKvoeV42YlqyW6NViv3HhjAeDPzGjMlMn0hj74WSgD7PbVMOSNcnPigRfEeZ79BSIYQXoAdIBK5wwRcTgaQ3eEt4AemsxKwIzKzDh5ah7clD8nc/Fz5ugj3SYlljkWPd9t8iOemVIf1CID03dUAYcTiwa9R+9tJIscWh7jJNItYCfJKzpDpEk/kMy0gUT+Hv/VnmSh6bVg2PLcDHfuYx2aV0Ax5rimYzQVWcKea5Uqe6jKuQfAEYVQZ8nMB+684cuXKs3/Yx2/e651rKV24lzAm2fxBEfDkLUQJMyF6+ku2IR3E77zRHiHr/5TrkhoLssncinfhF9H1EhmA31EEeHTvgFXPJv5G87B9IR78HkEPJ732FHIrTkIQ5lBQQOm5YW7kaZCOs3/LCOXnSxL6mx6gHmR69KN3eYaPfcj3plxpIaZqxkrEFIIx2dVUP0FIx/K0R/g2fewBDRdPJsHl4Rm20XMhxOrCE5Si4loEIJQsxJ7kJ3oTtKu1KLPI7stUULYWZjMVBKtHoDyDVoLVMaeYE8CC0ku1fIV3hoBWM2MGDWR+RL/9hSJ0G9JnOLe0zEnGM+KdpmhFXM/1oF3WtfAWwQSsCaTOUPBPLM8Z6579rvfJF7hohgO4bZie+uApZhczOezS8JbwiGeZa6LDGiH870qSDwJWWgaJmhyyPJeEieyKdU61hPCFYC0TGmw7ai/GwqzgcO5w47DKSkKDhH1c6q7GC625X3NA+swKDPzDLBMGhoVux5zbWIQ/Cx4P8YpWv3eddn269X4YlsxEkqUsLM9p/frr/u9bnXnT7j/EvEwE9TrLDpNE2l3qPUBNyMg955+CzfWcWp7OIKfHNJ7WvzxbhB7wJnAU1jT9m0/cPTBuNjJC9nHouJsOP/MuwEEo2k6X95LbWVknj/NQIQ7mxCg+FQAACAASURBVPi2p2Uh8YI5CWZCDpnasS3JTlO3XzbjeWLyPFPnNcR8A9Pz9wg7U7pPWsCj6My0g9MZmE6ft8CaPUX2sNaajLeAbs8XAmh+tOYnwu5fiY8k7sDv1Eywgq4mj6oChtJE0trYwJqqU8aKT7Xq7g0w2Ugp2MGxhAQDrOLz3ASJlB7vfpwNOMy1Zw2zkXYEjbkSWYgqMEriDAm2EskI1DXcsu5yeomzLhJc9socEyzY+IULYCk3qIU0sDP86zTi63i/IZGhUKq6BPkzI0uPBYlix+cjUVIqA7AJ12tov0DY0tzPdKBuGq9zDeXxhMhEKkosSaVkdKepqDFXNzhumASesR9nNq3FhRsv8l3XUzivYg6aVbOnmjMOH1XoIfP6au1yNAQzDK/X5htDoIShfQKy5mf9vc0dMJonB06VWtPB9JqmpEeG9umO7hFqRpq24Qieea91H3hdQz+Nkxtwo2TR6sBRzbL5Fc2j8Amh13Kv2o1eKnhhLoILi5h/3mrSC5c4uENpO5MMYCgsdTZISRSInTZVIoZWHwgSzIoNa33gfi6dXnMKM+hDiCXOHATo/IRYRPm5axqtSosScliTKV0Wg2O/VjUxWkMc3OK7rMMIDS+QiQ2BBhMHdiTcmencHjBSmQTmuoWNizUAqa4uk+BpAhDGw0zVHrulsNK/eV9tnuXE6Qtzs3zl2KNF7T2+FUwHKkCZtE8wxHj4JWXJwAvQZVKHlvyEh/Hekrn05prsrDcDJ3z4TEeOKNWh55NRPZtUmLO2MKNpQ6It/evgQKoYsX/hbvjKVkEdtMYPZAd1CKIqIDOYUYYh6V51K2uSspTuPZxVqlgP3hyr1dzmaa6IWxPTveYQT269xFX6kKNfQnE0q4NOLIL+N+1XxPNsmc957JQrjVOgpBik4PrWxOk1Sxa/AST+LtMa5uhYm+kEcYi1Pc60JTPbYZn/A951E6yYLKgJLCGpEIN4A2qARsnChKxTKnBcwW7eCQec12ymqmvwjqcWMucCcba+K2Yk3ajaSp0XbKM/66HuprQcWKYGqVUMHoLRGob/bmp41ISWwiTXe7VmUFBh3RKuUsuZ3AVqHQoD5xr6L+1akRczAzo2QXoKnL3GYVrs/n34RwYnRtteg3trCjXT1ydBTMTgiQwTPpMOvW6lJ6xLjXt8DythTlP40rq5n/saAjtsvoGxkKQKVsFDAygfsG01QC3lykjAmgzQ7gXgrs69HeXB1/gl4KQUoDpff0ZTY9uiTMhxaBO27Sci523YQkp+RlXvVEkJqD1mkXtiLCGS0+F5gOsJhoZZRm2eYWgfiiWIP6Nv5+GDUZj54TGxmjBH22nYma1hpI81Me4BOiOPUzH+DXjqyZgwtP8ipKC2kQlZw6yUAATDhio7GQXVI0W5Igx4MI2En+Epdl701WQofmHtKaMfvFIbA9UG0Vm5sfd1jPcM84Rl3rhDDYbp+gSJNZIS3DJc2UPZwWy8ibYQTJTkyMPkhJfkgUjydkWwzJC4GiMjdfZfDj2u3dcXEsEpjfhyCYnQANwNvPSiO88BTxxNPDt+iPgw8QxAV6qMIsJIJKHKOMeTpfBaQ2o28WwlEosohpmsKJrTbhcyS9Qm1LKHORxLZpJEhNApkogWJW3HtxmOLjrJKhOQEr0GLms5KUcwDOZzhPOCIAmLlaoz4CsZJsex2C8jksqO8axFiZlgT+uBjATAf6fpSVisSEfGCI84L2kosMS2o9ywaY23YWecPCVrSl/K+Xag+1wFtXQw6xz4HWIeyNy71hUtB8ngt9Zfb8Au8DCd1WUNjM+96YAl7K3VeLytKbgXa/OzrvHN7TRNRvBII45CtGM8APejpV0Q8Bru5MSeh5xiwJo4f7Q8E0La02r1uuP4ba6ww7CjJiJ8EdlwWhaniVu6M7QJvAkv6yVcrEW/Sxn51gVefFM0e6ZPJrUiSa/BCEm6SSpaVdMVqZla73X2vPg3ppnKbOlqWLopCdB9Evt+llrRgOaIAhnN23EV8f9VcQenIR2G3ajqJkx1Fy+PrIiRmMgo6OuGx/4ooiVm6Ox7knvhaGKqxJ2a27oWv4sENbT2sNYN2K8nhTvNCROh1OI86znbhFuvJ3HS2p7fdR0IBpeuUMtNB88OTuDZRLpIgKPiK1iwFq4izVgrW3OlxLXeOXqbKuWcI0slcFSH8FCNlZjkNYxreX4K02VDaAlXiKs3rwtLjXsr4EbGyeuhDk1BTq+d6i+wwYt3WZW4pedYhZ0019r6rGoPsTz6k2oWsycteC2aHEbeJixK6g5X9XiPkGyWblcNY4l+m2zxbn1hCCkcZ8+3th9IVpRqJD2rxanKK1lGMKDJlZoFQ5zk6HSWmsHS6XXp6oDUhsaO3Q9cq5RVeFRhgoiVoWRqRyO5UtXUTjJnxWvbA6v229g05Hp31OO4qDAlFJFt42A25ZmJcy6m83N74JFaDJsEE8E7ka41Tycv9Y1jmPNDARvMqIxQ6GgFvf/HMLczXN2FgVnk6PwicBdlM6cn7RBpFcY3wCehqITOvDjvhVVmFjRj6OchFBhxvDTmfMM1DB5SkBfbJQQMV83FQrVwjdDuAvPIuxEMpTNPD85yX8Y1yCW8twgaQhxk5eJV1hq20gAwi1xc3ZYSgMhgp11rHGYUYkRjRy1dShOECtIwGU3GnEm44/ijmjhE66jyYxiMzZAKzYKxf0NjiLG6l+HOCkTK9u2n5UQmTJYRW1f18ZDZh0C+F+qDp6nCZrRCRDrcatoaMoSN0r/OkAw/zex1PTM7IJ6PXhMiODKIDom6X0cd+2nimG7ri2q9NQRVPfNW76hWdgiesAyVnBGYEGASIMPIUlLn+o48DjEbrpcmXEm4eAWJf1wk4ToM1wqh4cffs+CQZ2y2CaZe85RddzRh0IHhFpO5xXkRhhcK9gfWsebxa6EAXN1LdLp7n0V8CcNC4aUvRr69LaeCt2rBdjHVm+tA7ptUl2xD1m91jN8hzku59G2WBBKQ19TCVVS1GPkIJYraR9G0sH3Y37RpcF2TUcobwCpsfdxCTth+N3JxpFb1mxDvUNamjnaj1l2p10YwwrCQzCNVTTLSjprwwpx9wnDBMER59HUndwC7UY9IEZ5eU5V4jcYmM4ut4bWmzAsx/FSkh/L6jr1cY4pxTq4DJo7oSco901QzDJpR3XAH2yOmdsdcFiK9z8trp/+BMMTi+tvvplb+i9rT0rWaGPPYRXJLsJ5NdGuDMIPkT5szPPtm2pHNs6TvI6+V4A+b/IpJpb8LZViBmdJhcgmGayBzB6/dlJb3hIuzI25u3r9OGA6DVjFcPVDrhns35ohbrUIz0E9qCJNebJ9RS+mOVNzCPizovgqRJtW07WKdce4Q2d0JO9Tl9YDs49o+1PSAUy071rnjudR2bGrZQYihdUtc+w3I1iiRQhoOqrk71zZyc945Ipouyb2tIT109+m1/HWBHZ0wUrcgtZISt7R4WGrV/N9oZbI/96i7KUkahlLOZu1LMEvpSqHQXc4aaRd4GXIjXMD7CLm2FOMkvOWrYfgCVgtXWfM4YbWgHACFnWfsYQRpgi3iskxYbjBgCGquiLPJH59XCS9IL6PNHZqGfz9qOrQmhzCpCZyEn9mlucOQ+MccDwmdqhd1+OqzNz1nhbcvH+dZb4HGMLSPhPu6j0LrjQYQqY7pwOo5HdhMIyMGBtpI6iGgEhGTk56py3I4YcnhgkVuu4CJQXsNOOcamzMjEP1cqNw6hJJPwnuPEctcnQfErDitkRLUkObL8/nWs8/w4trIAHUOx94COWrGO/xD+RNRB01HpxXspMwIhxDGyGxEjsZGB8GSNxuhxfepPNctH4z17tAMRD7idb1/ffHGvCexkP1SuITuX6MZH8lWJYyswuRnkBxHJNBnEQ7gIkwBuMqV8+eaKCMKWQJvePr8G/fybDfSNC/hjMc3BIx/RKa1lgNNXnTjSgVeCDxnktYpVDEaK9dmnL7LoTm+h25OamQVY6iaLl4jcWYTVGedRZjHSURa6hNhSX4eFucQ5s2GSdTCAZyMySqjefAKQOZejIUzXTiCDFATsNc2411zACrh5+d0mEYnqrfC0Ieo+hEiyltgaESJPYmJ5f7MkA7N42ACDw+7+uSopSUJHppWIkv8iEiqz7GjSnUioKQxvf2pGi+1SyQMqgru1cl5Mt8jw6OzRml5EUkTTh3sTWsrwkzZwCSexI0Kk8WwcfMnLjALBBufWqisPLoTx736we0k2GgdgBAKouEUPGUYzpobhlvEDpzamWAggWMT1gJ8xpK/aYT5UnfvHjwr+4qTaXvNf3VUglECYGkx+juSsBbtazkRZ2SpdAt2lIXnfC2Vlru0+QQ8bb12uFo9VI59Sq5C7GvuaqitpU3gMPLpeeqck7nzE0Eph2Nb87EHpWofc1kNNlwVhRAMTauEabZ1e9Ziet5La+8xX8bDHluYqAUzOhukW1+duDDjxLoOoswzF7ytznJ8EgNh2Lg5qeYi4IWVcx9zZPUwfRE+ErG3YGrLnxJ9wNqjN7U4LbTPUXkJfJl7LA8+cJBcU+uCBVUDpwAqw1e4KVY4LFo+DtPHoQ2ADM4VoVdoaYRhvuNyCoavEzJRQv/Uto/rThiiplqM6v7R8VeIaa7jlN5A/yM5ZD6PVNuekBfthN0EIKszT2RhlagXXZh0X9nFVHVPNUtOtHkmbWjuPBnglcgIOkzXqNJJaSTSQbanC4UYz1ZhV9XxfRK64CAk7rlTS2gGASETj1eX90hVvokBZz1MmnTCVgqERKd1jzL5mWdCn4XOj2GW65m5acI9Euoi4SvT7IqfFAZOpXNeDKHD5/7/D8PSuJbba/YYLRBiPYsFf6bwJ+Zxw5Z/aGbMmCfIkFMCz0mte0QUB5MXq2jtgKeDkn6tHCs7qOn3gVVIDuCA4SPwnZ211hMMgawaPhPWjGvSKgc+h6N/dbTrnlLKh8WFOebbs3bfCtv6JB6DuOcaSSl1fFQeIVrpmTP6MOeIB5hs1c5TdyayRI64fozdcI1CrZB4BEa9wbmHY6ekCS6rexkA0NnLG6QM7Arm1p+nKWBTC4omBV+GfQ6URpb4hy2pECgMWyoq0qQKumy4RcdEB8ezXs16G6KzxnIyXinE7PWTyZ76nPMAsgjqVJf7lDthiNmSJMKGITUnSW+Q+SLWwfdOzYiQbqkd9RNc4aFdGv8Mw2iaLBNn8ITFlcM0WE9RIszAk6JQJX47ZM37ZRpB+PwSrK2pkgnRNEXQGrWxpMmlOhGAiXLEC8DRyFlX5ZuEk6CHBd6SZyFNGGJVF5K5J8MLFvrGapeaOwuy1Ivg1lOI8zKXYWPhFQSanY1d7Ohk16ENqn4MkTYSPMgxyVxnDFZMDmmDt4GRy7hmAOHotHyTjTjESeTu77b+FfFr5x0xKjpbq4nsUpKPuzOf6eGIsbm+PVOmdjbINkzudtl2PZq0iJGbIKnWNggYnmQK0lINwfCMU93V/pcEWKqxALouBqFlVc7dPglqZSa8DEHPWWdqO6Nf4Dhb+8+Q55J2QcFix/jJtDB4VcLduihht9f25B/QdZLak3uM9s/D8CKcBoYAplv8ivN1iNW8gRrFzfgWTJLCkUSraAhhGbi4MzImYWttr4oRKT5yBgQocFVyAPu4gOqGUoLh7ntyNRdwv6ojtO29jF4Dw9Z0ldmoOwxv7eFWVr2W7FNyTFhMQyW5Ox1+dlLOqkzQGIAWCZRMwNGZBCyvDCTQ3NdRAS8TQvHzK4Wkbc5x2FFVbcY2SFQxUi3ZjTTTdpE8ltaj+oGFeYZ+DEvSQ9OpwsFwhnJ4YS/Ph4SR9TYYR1e2B3TFLJkbZbR9Py09LsMwErPeDDsaYW1aGYZmHn7tCjzhhzUwXLhEhIza9PgTMStAfqvR5khwzq5dp+RM3AsCNfOBCLIJjJGmwUjCUO+kTA5zWq0Ex/FdZEZD8BU3zydzO2AYmtjslXvIGhA6wkN8Cg/VfqAc+aIALjywBEOnuxuXmu4uohpNo4ql1oROj7ivOH4gRXKfkSY2Lxwmc98EwO3hRm2S9lVwnfxEVsaDq0BevYAFyUb8dtrVppo8eQ5Hq7xlgSlCyKQWRnJckZnhU8aYzT8YfqPqn151Igi92OPr4FpCT3beQ0LXN69fo82RAVob6t9tZ5JISvOZcQyyb0qozi1gb80+fcJtIDGmChudSAonUVUzmQ1rGGT/uYbse8r/LHhWvJMkU9Bt7/C7hJn7heR6AI5w9DMJZ/SZjt3h2k2CAzXLGlwMvB7ClhFLjYcMSqykn7iqJASIaz4fM6k+6zu618kd0F5b82GdUcPQYX4SqZ4/Qt1RxjCOa0aebBLDzX6Il8JAwmoLZyu18HrAmdU9xn1jt5eT5ojsf445B0G7CFNY86RmUlIssPR3JIaY0QAEBozvPphmsTRr4vZxmTtVWPN5PxOALYCO1jZlyDhKW7C3H7EGS0KtUdcGQLCgeolFrjtaE5E5tBMRSUg2EZO10yG809wxghsx256/aX2M0vT0yxJDIeBLa1cRVAzJy5sahKONHYVRiBLy61gHzqd0vkBKKmpgZJ6GLU0LS1riHaQlOAQLMwr+zHMnDIEjMqW1UGqs0WzI0DnYimzgzJxd8X7DJoutOmOTp3aNKfJc+5Ln6cxWSeyAYZ/nNftaYBtEpnHzLCsCCyhri9amG7g05YRXRsHZ+4rfCUPjoE87+qaMaXPvuZjYsgE8whFmiaAS2shcNEEEh150FIUE0oYeqLr5fVA6UP3lgYQNiJQuZzk3523iZO3GDoBZSpsr0wfx7M9gD44B+gnh4bTBFVDYNJdo+qTTVdl4BFMhicRx/ZJEYAWiNAcAR53E+IbYDcpSmGoxtTbCbQeCcZAHup0dJQ6Jk1JqdnfgBBGTCXWeywNDOOE6FO/Tnc07/X5LK+D9ujUwmCJAsLeEtQ0JLq1nxbyjm0i72VrbkdxFbQGudRFs0UVW6rY1+MVU6P0MEzaxkdZDpkHtN7qqxVrNWJhJzLPgmZbWnG5lHPi53sSRJxjK3J9nTnq2UbWP86LPgoaJ93y3LItQYMHcLrQYcl+W5DKk0gPS3Fg4G8qQc/ezkjSwU5MSqOe2xO+Jt8cLaS0uKO2AIaUIncqZB3He/tz5+pmIslaWczfsr0EoR6VJLvMXHY4aa2sttqON6za/3I6NN3irTG18IQeRxK7b7ElJ4JDyNVcu2kb1intPdsIe570aWSENj4T0ZFPrrYHc+JQM7z7n7IuggjGdE0PxPVabQ5ADez6d6YwPTktOLbUFmZy8tNXxjIenA9rrIP2l5jNhz8qdl/ZSg5eEEfcuPKbfa7Ew8dQmUmO7cBfuNZDIxFIgUysdmoHD7G+HIeETKgTbKVZoQGh8lLkfjnI8wbDQhlQjZm0Dhh7VaFp7qNaS5kULYZ6LGLg+MyMoAFfZJjxUpEQqEsBoN87RsTp8ZDtSJM6YixunH2bWK2cpzHUPYqoSgGsYRKrCDIGRPx+r4joH4TIxDcg5+IntTzrUDK855GCOfbBmcTYZjqXYvwMHGJfgY8QOjVYwdHRghbZC4WDHKLDAHBARSsLwKPwyDL3qYKBEypJokeR2NGQJDBIKz2dQQdDc2CKuWr5erMPgWPH8GichliOBNh3IpCuhMDA88ZmCrsDIn3NwjnZ968LG6+OsDa+EFv6E7619nzAMR7Zw0bjnd2bggdEp/KjFbI17B0qIkZmEo9DMRrI1O02NEgCs4pN7exF0oFEtZlFYL579HAiQ8JcrwhFpypI2oVaKObnstocKFdlCqjUZqvJYqpw804kpXY0IQOnZg4ALI70cErTmlDAsYZMdyr1nRx4a/iWmawbCPbU5dNPn6Q/ieCBC1HYX7/mUlcLJJXRix2ezryo5ByUZRgrnuUtqqVCPWsAJ27PxDadrpDyLuApnZiHBl87jGmmeMPTnmebMxbCozGo6BMPmlZzXRYSLTmJJd4ZjT3gBEQDw5lHrARTTrgmHhotN5pcDhrxS1OYLwZ/nHbjyJ8LwAPTghdf3bK6dMCzjRBXuux7doUgqStbbh71aHLD7WTCUp1LrdMAE8q0oHKsq7DmsikOy8O7j0/0i9Rr0nQDLFXUggVICXkHIQEdTBjjLh9T41wdEH0WXwnABO/b5TKgb11WaE2gVrqtt6SvgYduEsI+nFLZi5WerqY/R7AjD9KTwvCVWQbvYzCI9/2SjW0jXnbTK66jd8fS3EMs5rRmYwueRxs69qcR+mGT2hhgcm+8MA/UHwRIM1p56EYX2gFpmvoSCnKdaiVXrwR6dqwnT5f+284nfPCNq1+kr6+93RJ0E83X6vLqfScNp8/Z6bDzq9ezZ8HQV6ghbMaZ6esY+i4Ydn1nIBkN/EgwBKBkuhWsHIUZrqvPc+UzVA5fkWTOiqTq9CRA+DCrip8ee9hTK7y1ABMKEldMupsr3CFVHVK8fe7Ttd3A4x56CM4REFZgRA4LjCkYTfoI4qFYJY5Wpxj3lFjCttrWfaQ1Y/eTFcFvZ5DKRR2Mf/Tv+oep1LmZPSmUkU/F1DDQPVAsqjWYFDFdInSU4nmhAJMloFkYYnzUyzBhsiW5txhpgjB91G89z5jw2W26ed/w26ygHcBTKCjexJvpCqK1haFfLeOhzNc5mgZZhaBznHijkmHHL7x64jhyMOua5BCaUo15IM2fWzXnegGEpDjgw919mkgvqlVHEkhsupPCguWLTq5DzkulsjSlteK4B9VYKzA8VktPm1WBG1ThcHnSk7xacTJUHx9BYSGyPNepTSDh+xlJ2edGlDhlgcuQFAlO1a0w4zYVEdhT38qxKOgKTvoEegwRhQ63nSxheWuOwgoCeR1Myk5BUQ4KLS+erFhywtP3Kvbq1Wr9G2Dm/wuNxzlBbA4bUUU7GnIwfsZY64GSQpisYSEyyEDr3sPI/MYIrxiHsS597Pxwv1xu4Rm1CeIfjfRB3ylqFzOyiRmqzzYJnG7/kH/PfeIKh4ZgwTOyo498DB/n/R1Gd95z0lbB8pmbhf/GznNPj6bwLuDMlWN7wWJYWSW44mY1sT6vsxghLHmHQmSoTl9j8V4RFAqAduAI8ZDAgwEtmBDmrnhsu7+KkOdKaDMpBkrWeuSm7XD0hLrw3ApMJYEswsVe/BoaluS0JmgBZPHZm0HWhVoaLr2Pt9p0ACAcnD9aSunTAxwmGBzRbtCnlGTQDifgYx6KjVPSUtxQtRZ9S3gfEhWxENSX+6KvSWXkPp8xMhszP5Mk/YDhSEJjIA9P5TukKEfA5i52DS4+XVg6dQ8LQEv9JExWD4DQ+rRqtw42M6YTO/h4s9SeOFRjLPnEKk2xVoY1bYBKmJzpkJqi1kmQ4vc7SWp75wfQW29ibE69BCuemCzVT2s+3V5YmA3KGdfzc1Xa7MGP6dqpiPb4cZ5An3iFZH2/mZBz9HiXZlqUAY9jyDJOJjwSe/y5qIariJCpknknvgQdbnGdxra/AgjeI6Voqx/GjdKMbM/AKF+6CrWFTQkAhNn0tR+7FI2AYeRUUHeW7PQlDiPDZ8WlUVL1q5tNndDtgSJjT97SmrZvQasascfoaxXvso/dE0QFJ6f0Se3h2Uq4DrgcMebUCws1epb3b+c21BzugAx5QJMff+UzEEgP3FF3jOcAOzX6/83PsYxt3rHDDJpEKDMV2KQDM1OjDkKla9Hsg1runkc8yrsICotfgd4h7ujNlPqe53X6ulw6dLqyIb1+z2eQ6RILw1srJRJliu8eb9aFTJ7lGUh1SsgDltq9+S3eG1gZWqqETCpQ3+km94iqKRdL+/Ci+IiNUFhLxYwETH0+u7x6VzhloZJy+pLhwOjhPnwAR9jpgSGZxzRIShq318KeZ1YXccSIwYUFfDQoKtXJvVu+hUToj0cTrKA0R9C1Zmlq7zzgl9TV9WausaUrkUFsZLOm+SA+tjRdn83mF2UPwXPAzPAFiTa9kh719C2Zx4gv3X4Nv7Hi9gmi1txEENn2IZ2uwIyU0f3/WohOG1L4ShvYRuibk1HTyWcFgLSVicS4lQ2NN06qNhXvgTSfmeW2e4Ro4r9CeN666LyDSe4egjqpAIzqdhX0Qs/mQvo2I5N4nszExE7mXEr+sKwUnVfIIgUopS43Dek+GmHQr96GGEvBkKpfQ0BEKz70mKcqOTjKp0ILASEtZJFciUzIvw8AwtObkcmXDcMHt6w1dqu10tC6lkesnVGb/zjXTK369sbL+30uaDAnIGsPld+stn0XGKs/MzrswUwvNMMrndyBsGVfW4u8OJdtstAiidtOS8IFUsZ0rEUmC4D2vY4rVhpyiC3B0jNpZaW38263yrIUp4a5OmOb8YpR1Nvnl1YabOSCMHmmPPktRpRgJvWPzTc7/FOUEmfnAyY2zIdyE5nWi28K17jXq85UVhwrPGSAFhp66XbvtVxYg2Z512NHqXc9Kp1HNjoJAQcYBZaE1IwiNIKS1QpwzQErrOY1TC0q1MdRO9mJM6tllUykZWZeMz50qMndedN9C7r1iDv8QPg+eKJ7TswtL+GfZShX5dD5iDvKqmwiP+1z9gmYWAdK3chAEGYRToIkkb4chmSvVc5b725Fns8XMtpd0i/Z5hPADbNh7hMA3EXXFOHEnytpaQ7bYk4BYlMzEZ0tkFV3RaSnnvLOMBTWGToO1GXRjLvKsi20GuQme1zyrV3d8X9joqzndbSzp8PnnAsJhvWc/jHJVnH2a5abluNz8uIfnGmZ55qtgHMJ3vpQSKW3BQ8VnuEeah1U1w+b8TAdNblfCE39fW6YPsA5ES8cR6yKIqFhGwvZNlA72rPQsdO+L527R5uCQRKMmkkgeDkfOM/zc0Y8YlmHlvBB4jpX7NwwZ6w64yctuycE9tTbRxHE4DmX7A94/129Flo1bztBwzKOxoxeJogVbcOa4ZkLPZsmpnYqZHREXYtduOdJjrQAAC+tJREFUmFXizRUMJWHIZ0jgDTtLYuoa7S/RswELmRFKi+5xjyiQxmi5n/BqcyWcszqDYAD0Iel4QpgdPxEUruNjf463vZMm6Th3w9fj948hBfH0lVhjpSwIZ2rgIq++cmt+tVQrTeAkm2m+sVjiPZyZSUp0tIFOKKvijGJwQ9QaqA4RiU5paBWc//KgqRGGOmJJVSLvkEyw8yqIMzWLBFCXZJt3cw883C4wKr2Lmu/p+FRSU66hwMYta0UvheWio0saVsX7hI3hKjSqlLpJiIMITGwSzKl9BJHw/dH+DIdz/YIzzHhFuvqlicxM2Qjv46r4rPrlbDWwFphc5eSkZASSNNpnDU66SMvwsp0ecy5Ym6g+Yy9tBZGk5tU46YY48w01NWlerVmROYqSjmcCj0mookHiD/d6avn9bDCiJGy+k7zn0Cwu+TB67WYMTTuhBIR2UvXAvTshVUw04DwSNYjU8MvD2S35MZ12+B2EfJhUWnff8ubOQi+ug6vgBolUHPRxIECvdUrLiybBzQdIgJG7C6kHeKiQ9ARkKVSaKbQtB7feP1PXuXZrP0byIfq4PTtNKJoOlT026NEeZq6eESu1md6j5Kb21WwgzzE1G7IPSxQi5PK5zr4ywlLb2puEDCq0gkIVHaBjK0cVrdX80VwocHiOh/PU+Ebonz/WppjGv/qPWYfhw6cpbMwqT76wiLPCUc9zaslewwAep7Q23omvzLP2x2mCoCf6POZZMmoJwwwshIHDSBnTE6ZHjOk3NWr6+QK+a4RzmEGpUS4s3G+4+vYqgk6AGASU83BpE6nKpJK04tm+P9Gb7yk2LNXHJKCDbrj7YE+MavuyN/IQwKSpJPeOzMBO2lrSjFjy7HNzDoX9ANRejBxXSNF0nF3VziGppOHo9KbW8ZuKjfS/GyZYh4AvzL2oaQIMZk/wTYySWpqPsDQnLXStRKExwtCY75AsNbpuq7dq4bh1LpDZvSBK4/X1lpAErtpgDiKLki7cW3ura7DBjCp/zNRm79kM2qIT1AzegCFK+SX0bZAxSkuZRi+HgzbOhONTs4B8WhSmbGfHnhk9vs1HEqQFEg+sGXoINVAwN24w0sN9pUsg8zpLMLyBxWtHsaXeC3omTDkAhWBoXWR6ux64p8mRw542JQmTG7PUZJ6FF701xnHsclIMx5Q6u/SdU50tsdvxw/yG5JA86P78GoZhDTLz7SHAGLQknjmEBSOQ/B37OI4B29BKYeOl96s98blktDOT8iBgDWckBa90NAz204kQTlvIxHFEtAIzbW7rDzYzMv/jMDRh7WqOKZjOQTQHgRKGfoeaIns5StrzeZqp41jbYO7IMm5xTvh/1rAYqgFpejUMbzpnN9Gx8cC9iDiCufTy9rlPMalWwdNUO3BEKy2dT0aoDub35M87WCH3GTAkbq/nZweOaQEYhnMzHmljefzWbO3A5d/GQ6am93gLq+tzBkR3bsKcqUN2QiARc0++INqAWrvrUI5jJip5nFk0JWFmK/L7a92w5xmshauYrFKUPSBRO77ObETEGtbTGvI7rpIFSHaG8VuuqSFj/4LVv3NPMhsEww2Hy+KwxMnJuX0Yz+tMmDaq3LDCtraOl/asyDuQwbB+iLCyZT6lWDgR64SFIfkMVzN4M40lZtXhwMgcTRUof2grV66JWqVbInIcMWRQ2vuvhMUzVvrM1jHW83taFoh/lMajVR5hWvvFmHXD5LOT6c9aw1nab1trtS/hec+GiGHtPST8j4jQ+N+8IbbPowDqj4/2i5ptidYXFi7eGu5+AGvsv+GQOh8rs6ezCdqg1bdWk8QUimS+sMCWeWvUpYwRW8tAfG/Ehca5eCBI1XVNjkJoDCQUFe4EOBgJOYBuwid3bngg3o91huTL+hPCAMX1k2MboU9G3HORYMkQnPvw3C6v+0w4t59Mw1I3Ycy1ngz+JqJ5zolJFusxpCfp3yvt3IGdOo7RxqbCUDm+//a/gW+cQ7hIuENM25MmDJ8jFLHexBPh0U14BP4N44U1p4ThLX5nRGy9ASOu3cz3inP1GnkfTsW+a/ChuF/68sq0dbDbwwTGYbYIf7WPejJRKFo4R7oahOd1v+g0E9Cp2jKTrD9npl/a+VSPjPReDB1+Swv3u0olFwOqWDSRdMfvdOz497aN3Tvh2Ngb9jgvsVkxg/cUIIz1e38A/REnM2mQMeGFzq2l39d8Lzv58MUcBzGfULIQGNW+n8Wzcb5DBRzOcF9KZK4CAfc0z9hDobROPicMoYNOjs08ZUtIJwJFLw8yednnsdmEXRC7AyMJh3yvjjGNfwnDEJHhFBQe1gbUAZvhUXqCOJdxyVpSaxMJw60Gz9UwAqCbyHW+PHuOBe3ZWvcCr7ZgaYG01XDS96/2YTi/J9MMtuAgmAskSeve6/Iu9G4qBVW17hsPXJNbzkUTEXtMJThPb4RZrCY6lWcen7gUSWIy1hjimhHFxSQrlg+7/Q+2rSoOhgd1re7cLNVrEQmvmKPfuA7anF0mQwEMnBn/sP6V4eZxm6DMGAkTETNq5g3OLTglkVd+hWSUu6i3sS5mvNfM8U+tSYxl3mc0hX0ly7MtMNU6U4vdG4JyUpc8jXRkQ+Yk4H6atRkvY3rUXI0QeytmhhKm099k9rJUSxL9KAlTOhGDwEpw7LPbwejsg4pnhANuqpS4mtjBc2eX8T0Nak4Ycn2xT/pMoiuWTV3jh3+PsOasc8caqVSsWK8zLzd4H0oL6BewHqhT2LmupGf2qk3DJrXDt+HhxtXK7G2U2muO6QqvtRExFa2s7Vwx7PP/4+l7HsqKccleCJn1tmcPqez3KhxoqeGsAaRVMb9PFPM63/wPleoyNQ3vmtWiVMWpjtKk4r82E3IewtBeGMSavMZYQ+7xQO4nWEvC5t9MISYzeD6bJLD8PM/VpkmS6YkXqd4bhjxXVAV8YBgJYtnV/TiNN2BHWOQZnnvLtQ++Vpy/0OHcT77jv2Pst8CQxHjiNE5crJTgbLJj2J844sYG/izP5tJT10T/EobXAdmk5zBmI9qR9PwGvQZjvoMqaAB4U9UqAskZm81Nz0Ip858MRYoX4pR4JG4D3FoK4Etj+ZIdlxmK47cq+cWcJNaEauvww5DAkpeSm+dPquCWQrMi5SI015c6n8Q2DsUaB2cjyhZ8KvapC3UP1IsEKO1yDixj3wPPfDLPQhc0L9rhhmEPZXl4IIm4NGF2Otn6EavZKeVd7/mABMCxxgWmtK95zjC0ev+Mb4dkPHCrcDiRA4bnT5jP0iQddo8Thhnw6sjBnJEvk0oYGpvehCEEP78X5wMzIEd2eP4R1o315F4qxvBJPvBMly7F67UY9vutmdhJvz7bdszfAedU+mGrTw20BWb+reO5WVK1uuvoxELVa21Um57n/N6e2pJU47ZsSvYh1AnIYWZVkY1HmjlMAVaxUCiBtsL2C+RaJ6JRRRRjInDzVjZFX5hcxH2t2TLf8ZiNXFf8bp5NImoYMo3X8XyipCTUICr9Lg2eJfgm8+f1AvTxkDhYD7TrGVFvJwKffEJeejJl1aIsIBlvDRzYS6ThsfUZ9ygmPDBxHsUwjQw3rn5nFy8EXicMZ7EsEuvIGpn2+AIiWY+e/vgfUKKk014wBKNXJdi6rJumshmecDVzU5ZxjFPStMk+E8LaAtRCT8wNYCfu7FNRgqH9YWI8MlXX0NwJQ+Ms8XDpjMi073W9/id1/+i/SA5Ww+mVNosLiHZdJFXbr31k5HeDpk/WI/tSBrPoQB4QnJKc0zar+f4Gy7TthuLzF2vv4ZQlObAE/LgnYtbYwEzZR6R7YOO1JVvVWuuWCc4Dwi79PcflfC8BQ45r5S4dXmRA+y1785kQJlfMlmNUwCdKmLXbDvux9sVdMVa8K/kYu3Q/DKcdp3xPDa0GHo+B4eSiaBUXThgizi/zELgnJ4pRGV/w6QUbfQOG9EIZhg/UlLczW/VwRAYUOzx6B/N8MnNy42U0jSMoGesgHpvpdvGWo4KHtqNdcEy3R2BrxfSL9N+vYX8CZp3c2+snPKRF0OdXeI2+iKuT0d7EQ67dLKfWR//0PwK5GG0E0c44NQAAAABJRU5ErkJggg=="},{"background-color":"linear-gradient(to bottom, #f4f4f4 0%, #f4f4f4 100%)", "background-pattern":"" , "items": [ {"x": -214,"y": 97,"w": 878,"h": 212,"type":"text","text": "Page Title","font": "raleway","color": "#a10705","font-size": 28, "font-style":"regular", "justification": 0 }, {"x": 1534,"y": -153,"w": 253,"h": 392,
            "type": "color",
            "background_color": "linear-gradient(to bottom, #ed5353 0%, #a10705 100%)"
         }, {"x": -209,"y": 333,"w": 1992,"h": 638,"type":"text","text": "Lorem ipsum dolor sit amet, consectetur adipiscing elit, sed do eiusmod tempor incididunt ut labore et dolore magna aliqua. Ut enim ad minim veniam, quis nostrud exercitation ullamco laboris nisi ut aliquip ex ea commodo consequat z","font": "open sans","color": "#666666","font-size": 16, "font-style":"light", "justification": 3 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOy9d5BkSXrY93umXnnXXe29nx7vZ9adwR15IgEiJPAoBE8AIxgkpCARogCSIHBQBIMKBkSApARCEEiJBGEIUAgRBHgCDjgHnNtxPabHtjdVXe27vDfPpP6onp7u6Z7dWTM707v1i5jY7Vf5Mr8073v5vvzyS+nLX/7y/3Dp0qWftdvtXurUqfNc2MNhW9Pv/Af/i8o/f+lyMf2FLxRfVP7vhWq1mrt169YvqZcuXfrZz3/+830vW6A6dQ4TJZ+Ptd+2Xlj+7V1drhNvveV6YQW8N0LAz6r1GUWdOu8dIQSW9eKUhRDiheX9frDb7V71ZQtRp85h5UUqC+sVUxYAdWVRp877QAiBaX5yZhZQVxZ16rxvhHiRyuLF5f1+qSuLOnXeB7WZhflC83/VqCuLOnXeJ58kAyfUlUWdOu8LIcQL/gypK4s6dT421A2cderUeVdeuJ+FVVcWdep8bKjbLOrUqfOuvOiZhVVfOq1T5+NDfWZRp06dd+WTtjcEDouyEAbJsZt7rM+Sasd3/CSa2/7Ri2MZpO/dwSjpz0zjPnICpZqmXFTwDXQi7c+FwtwjJH8PrmbfixS3zgtBYFl1p6xXDyvP7S99Eeflz2OzywCYhTS5aJJzv/47hI73HPAwvkh5Kqz+/u+S38gBoG9GSC6kaHn9zE6Snv/x5+H+fyI85eO1f/73MFNRvvsjf4vXv/InOP0aQsDir/w89k/9zwz/t5c/SunrfAgIAdYLXLGoK4sPgqpx/Fd/g2DjtshCEP+Tf8+d/+nv89mv/r9ozo+uKpLq5vg/+9Wdv7Pf+m3Gfu02l37zV/corWrX38TzOWVHXiNfeJLHR6rd6nz41GcWhwdJovELP4rjF/81idlV2k71oKe2iH3vO+TCa9i7Bmj/r/4imsexc4tVzrP1Z18nM7+Ma+QUbT/wKRLf/C+4zn0Ob3sDAHpqk41vfoPCWgLPkVO0fOYtbE7b+xKxuhYmE7fjbnGz+G9/nWo6zvyv/St8x8/S88Of25deCIFVzLD1598ks7CCo3uIts//AHa/+/21UZ0XRm1m8cmyWcgvW4APhGxD1RSMShVjY5Kxn/hJMstpvMNDFB/8OVf++k9QKdTsClY+zu2/8d8w9e+/AqqNxDd/n5s/9XMs/8f/QG45AUBx6jpXf/Svk15K4e7uJP3dP+Tqj/9tionCO0nxTHJ3vkP0G9eQZBVXTzeSasPd24+ztenA9NW1GW586UdZvz2Pu7ub8tQNrn3px0iHt95f+9R5gdQMnC/qX90p60OmEnlINqUQ7O9AadC4/Du/i+qsGTzb/vJfRv/bf4Wlr91g+ItvsfRvfoGS6zSf+ne/iGJTEEKQ/u7v8/aXfo/2nwahZ7jzkz/F0C/+R9ovDiIBXT/yRdZ/55e4+09/ldd/+efe/6eDzUnrF/4itv/9N2n7wR/G6deAvYNBWFUmf/4f0vRjP8fQFz+DJEkg/iot3/497vyjf8IP/Kd/Xf90eYV48TOLup/F+8cyWf/P/w8ZzxMDZ+S3f4Oen/qnuEMuJASiFGf9z69TyRTRmtpxdLWTn48irCIrf/hNhv7vP0Ox1WwIkiQR+MxfJXTqnwNQGH+bgtRFaLCBajK5U2zwc1+k/G/+O4q5f4Db9/4+Rw7i6VmmsbXI1qMkr/2vx6mmUjvXXac/h231F0htlGloc1DnVaG+dPrqIgTF8Dyms6YsJJuDY//yN2i5fBqEIHvrG9z5J79G95f+Br6+HirrUWI3H+F881Og5yhlJDydgacylZCUWhNUUjEqy1Pc/fs/va9o98lLSLoJfHjK4ulZglmIU95a49GX/wGyvPdHbfg8lKtAXVm8KrzomUU9rN4HQVEZ+Jl//GQ15CnmfvkXGPjyb9H91kDtghDo0RskyyBpQbyddlITUXxvjTy5SVhYlTIA7p4BFG8L5379t7CpH/1839bQg7MpyLFf+jX8bfUYyq8+n7yweofbwLkLxeGgtLYGbEcxKiRY+9qV2o+SRv/f+nGm/5efp5h6fBSDIP7V3yI+XTNu2kcu03HUxsSv/V7tE0EIECbz/+xnWPyTGx+KjMKoYj0VXcmq1pSVHOig9wfPM/kv/0+sx4NQWKz+9v/GxL/7Lx9K+XU+PISo2RVe3L9XT1kcnpnFOyIx9A//MVf/5k+Tu/k5bJpJPrxG0+f+CtEr38G0fpzmv/aTDCwu873PfYbGS+exsjG0I5+i6WRHLQdZ4+Sv/iZ3/u5/z9tf+gbBkR5yD24id13m7E+f/8ASyp4G/B02rv3oF7G7JI7+8u/iGz3Jw3/xM6T+7AQnfuXfMvjlf0Hly3+P7/3Ij9J45iilhQmqNHHu//g7H7j8Oh8uodde479e33xh+Uvyq/cel772ta/F3nrrrdDLFuQdEQbJm7fxnr2EzfbsTwQjkyAzOY3sacA3OoxsVUhPhQmcPFazEQhBeTVCLrqGs3sQd3sj175wkYF//hVaz3TXirJMCvPTlGJpnN0DuDtbaisT74CR3CC7miN4YmiPU1ZlPUK5qO64e5u5JKlH09g7+vB0t4FRIX3/HkLzETh6BFmRQAhK0XnyK5toLZ34+nuQ5PoySJ2Xy5UrV+KHQ1l8YATLv/mvsJ36IVrPDu1czY9/gyt/55f4zLe/icP9MZlk1anzArhy5Ur8E/KESDR96rPc+rs/QaT/FP6BLsorc8RuTXHyV/6vuqKoU+c5+MQ8JY6B07z51W+QHr9FcTNJ4xuf4cQvnkJ1fHjLoXXqfJz5xCgLAMlmJ3jpTYIvW5A6dQ4hr57JtU6dOq8kdWVRp06d56KuLOrUqfNc1JVFnTp1nou6sqhTp85zUVcWderUeS7qyqJOnTrPRV1Z1KlT57k4FMrCqmRY3Uq/+IKESXRp9cWXs1NckfuTcwf8IHh47yEfJFqCsAyi0TWEZZAvlD9ATgdTKhbRX2A8h3dDCIt8vviM3wT5/PuLm/rM8owc96fCpLfWyBQPOC9GWESXVt41n+WlKK9geM3n4tAoi5WN1J5r5UKWxcVFcsXag5DL5cimYiyvbSEQpOObRKKrmJbArJbJ5rJEwotkC2WyqRjhpWWMfYO9trvT0qvkcjmikUU2E2kEYOoVlsKLLK9uYFoWmUyWWtgLQSabwdQrZLO1MjL5Erl0gvDS8oEPlFEtEQkvkkhnyReKgKCYTbG4GKZQrgJQyOWB2kO/Go2wuhlHCDCrZXL5PJFwmFJ1b97lYo7FxQU2YknEdm22lma4euMOa5vJvUIIQWJzjcVIlIph1qKNZTKsRiNsJTJUSnnCi2GKFX2PHJvxNJahc+f620xOz5E76MEBhDDZWF0msrSMYQn0SnG7zrV6lQp5stk0iwu1PgEo5lIsLiwSS2YQgF4pEg4vktn+XQiLzbVanrH1KG9fHWNlvdYupXyGxXCEUtUgn47x/e+9TWR5Hb1SIl+qbrd7kUKpSiGfI5tOsLSysScSqhAWW+sre8ZGtVwgvLhIOpsjXyiBAIFEIZcjl06wuBihVNF35SFIxtZZXAyTK5YRCIq5NIuLi6Ryxe1eEeSyWRKba9tlCUCQTcVYmJ9nfn6BXLFyYLu+TA6FsniacmaDa+NT+HxeHty6zla2zOStq8ytpPB6XKzMPSK8lcOp6Fy7dZ9yap1vfvs6bq+P69/5U2ZXkrhsBmN3Jp7K2WIluko1n+BPv/ZtNJePZHSKqcgmt69fw+b2IVtVqqbJw4np2i3CYmLiEdVsnG9++ypur4+b3/86k5Et3JrFzduP9sTbFMLg+9+7gsPtI74SIVfSyW1FufloEZ/Xza2rV8hVzZ28b169gqE4qabXuflghkpqg298+xpOjxdVebJ1XVg6N67fxOcPoFfKCGGxsryOy+nC4/ET9Hv21FRYFbIlC59TZuzWfQQW3/rjr4LdzfL0Lb4zNoHX5+bGtTGEsLhz4zqWzUVqZZq5tRROzUmouQWHXdnXP0II7o1dp2AquB029EqBK9du4fT4WJkZZ2E9zerkOGMPw/gDPu7cuEa5lGXszgT+gJ9yqYhZKXB9bByPz8+DsStkKib3b14np8u4HTbsLg9uh4eGgJdyeo2bD+bxe53cuHYdxenBaXPS1BigmFgjvFGblRZTq4TXk8zfu8nE4iY+794jFsxqkaIu4bYZ3Lw7haWXePvKGC6vj5WFOSqmRTa2QbZkMnvnGg8XN/F5nVy/coWSYbESXSO7Mc90NI3P66ZYLJHfWub2RBif34+wTFajK4Dgyje+xlbewG2zuHH7Hrn4CpPhGKFGPzOLS7jsr96epUOpLJYWFjl+5jShUBOnjw2wFFnDktycOj5MwOdmbmEeoRfZTGTIxOJYAvoGR2kKhWhtaaZ/eIiW9l5kPffMMvqHjtHaHGLk+GmSK2GamxtYXl7G4WvA8Yywe739tTLam5voHxmhua0b2cjvSWNkV3G2DNLaHGJ49AhOu8L8XJhzF88SamrmzHAbiyu1wW1VMhj2ID0dLfQNH6OaimEJQd/AKC1NIWy7lAWSQtDnZGVtk2BjI49DYGiaHbvDhdOh7ZFDoKJSYW0zQT6TBaClo5+OliY629vo7B8gFGrCp0lUSymWt5KkYhuUTZmt1U00zY7b7cGm7B9CQs9TwMFAdztNLa2U4ks099VkPnXxMqszM6A6OX7sKI2NIdqCTvI48NphbStBKBQivb5AtipYX13FRpWVlS3ylo3Bng6aWlrxOOzYHQ5cTjtzk49QNIXVtU0quRwVU8Fut+N2OQ/sJwsHJ46NEPR798QfkRQNSS+yEc+ST6cpJqI0dNfkPnZ8FHV3XBGbl5PHRgg1tdDX7GYzVfvscfpDmIU46UKVxqCf+flFzp4/TaixkQb/k3CJvlAnI/3dNLV1I4kylVIetz+A1xck4HWjHNCuL5tDuZHMpipU9do00dB1ZNWGrKo7QXDtLj/DI0ewKxJHj0pUEsvIypOo3vLjhO8Qukw3tqffwkRICn1HTtFZKfJofIz84Pld91pUK7Upo6xuv2UlGelxXz9VhiTJWObjqb2FZQlsqkzFsPAoMlXdQH2cj6xgWeZ2FmLn00Kx7X/rSJLMqQuvUcplGLt2jYtvvrb9w8H1nB6/hatzmCNHOkjGbj8lPyi7A/7ICsGmNkZHR2t/ygpTt29Rm5MLqtUqNs3+JAixJGOZNbklCRTVhlE2anU2qwhFRZIE8k40KAlklfOvvUE+neDK21c5PdJCR3cfo30twCgyOlc3lnby3I2i2ukbHKHZrTI6ehR1lzKXJGnnDA69XEbgRVLVJ2NgFw9ujtE8dIIjXXaS8bsgyzunjlmmucfWIEwDc7tdddPCtf1wa64gb771BrG1KNdv3cMnS7VPUXXvDExWle2ATLW/G1p7ePDdq0yUkoweP7lPtleBQ6Ms1lfCTChFkG309A5ze/wWmaZGEvEkpy5eZjrx2DApMdTbxd2792j0e7B7ArS9j7OT16LzTHogl9iid/gUM5MPMZAp6wLNZsOnGdx/+AhRyZN9D5+XircdOfd9Hk3qVAspZMnF4Ogo129co7kpSCye4fIbx7gXBdnmJahVufvgIVTzNHT0IEnGgflaZoWHDyZQNTtCfvIwqE43mfg0kRU3vZ2tO+kdDo3YxirZLZOC/s7H8Mman0aHxcPJaRyqRHNnH/6Ag6nJCY4MDfDg/gPeeuuNnbe0rLoIueDOvQc4VJm+4SEK8zd4WEmRS24xfOIyxaW9n4BGucC9yQVsmoqiagRa+5i9Psa0nkUSgoEjozR5ZG7fu49TVegbGqSY22BxqYHBY8e5evsW6eYQkqoxMjiAoWeYXYjQ2xEiMTXOZCXORnSB5uGDD3gCsNtVNtaWia/qVAS4GrspT11jwspRysXR1MYnbUKVB/fuE/LZieUlXgu6iALp2BqR9QQKBppmZ6i/g7Eb12kOBfE2tjyzbKNSpFw1KJdKLM7P4z15fO/M8RXgUETKEpZJsfTYoi/hdDoRlkG5UsVud6CqCrquo9ps2wNWoFerVHUDze5AlcG0QFWV7ZmIiiyBrhvYdr+lhUA3DMx8nImVEqMDLSiqht2mouu1/FSbhl2zISyTUqmMbNNQZFBl+UkZho6sPClDVW173oaWZVIulVE1O7L0RK5KVcfucKLKErphoNpsICzKpTLIKg67BsLEFBLqU9NUIQTVShnDtGp1VmQMw8RmU6hWKphCwumw70pvUS6VkBQNVZFQFAXDqLWHZRpYyKiKhKEbKKoNEJTLJSwh4XQ4kCRRux+D2fAWJ48N7ZOnUi7VynU6wLIol2t11mwqpmEgyQqyLNXaS1aoVsqYlqi1gVKbnZTLZSRlu+6wJ09Tr2KYAofDjmXWxoNq07bz16nqZi2dUWtbzW5HkmSwTBRV3RcuUVgWpXIJRdVQZAlFVRGmQalcqd2LhIQAWeHhzZv0nzyFIiwcTgeKVOszRZEpl8uAjMPpQJbY6VvN7gBhoaoqxk7/CgzD4NH4DfpOXsKrKWzM3qXoH2ao3feBnpsPk09QWL33RiW9yfR6hVOj3S9blDqvKI9u36H/1Blctg/HthCde8hKsoxTUyiVDc5cOI9TfXXsFp+gsHrvDXughVNPn0dUp84ujp8/96Hm1z10glf91fTqqK46deq80tSVRZ06dZ6Lw6kshMXM1ByWUSGeyCCESbly8CrBe2V5YYa88ewl1emZ6fecp2XqxOKpd0/4ATDKaeaWNvZcM019Z4n5I0MIYptb77QqvUMqHtvn4TozO41pGsRiez1Oy7kYkbXEc4pgUK688wrPTr7lCvtE3R5f+68LZqdm91//EKkcJM8rwqFRFnq1TDKZQjdMQJCIp7at1xXSa/PcnVh85h4IyzRIp5KkszksIRDCIptJkc0Xax0jBMV8jmQqTSaV4OnnSwiLbLqWPp6sDVjTqJJMJiluu2c/dQeVcpFkKo1hCRAWpVKlZqE3zJ37q7qJZeqkkkky2TyWEFTKZXKZNNl8EdOo/VauGjty5DJp0tnczvF2RrVCMpmkXC6QyjzZDyGEYHn6HjPhdYplHRAUclnSmVobWHqVcqV2b0U3KBVypNLZ2m+mQaVSIZVMki+WtwevoFSotZFp1fwrKpUKuUyaQmlvG5SK5e02qJDPZnbyBTD1KslkgkKpTKVUppaVIJdJk8nmSSSSCCEoba9+6ZUyiUSSYjFHOl+iUi7v1L1SLj9ps2yaVKZWTjI6yb3pZfLFveNBr5Rr/QFUy2X0apmbN8ZIJNNYezZsCBLxZK2O5WKtjbb7IBlPUtzdDtt9mUomKZYq22O1QqVcIpnK1FapykWSydQB2wtqK33pVJJCqYJlGtweGyOeSKIbL2/fzbNQfuzHfuwf9fT0uF62IO+EXkhy/c4jbCpMTM3R0dnB2vI67S1+5iNxXBRZyxg0hQK4nvJUBMHdsWtUhEo+k8YdaGT+wW0yZUFydZGccGGkl5mMbKIInYmJKfpGj+NUnjhuTYyPkSyZFNNbLKzGOdLXwbVrYyg2G+GZCWRvEz7nk3ILyXXuPFpERWdybonO1gZm51bwyHkiWZlmv4vMxjzLGYuliXFMRSOXyeANBvn2H30F2e1jIzLJg7l1XA6Vh4+m6evtYvr+beIFnVJ6i8hmjpaAnavXbqJqGkvzM5iOBrpaGnbkWJufoSi7afB72VqaYSmWo5KNsRIv4ilv8o3bC/icCrfHrlE0ZPR8nNVkFb+U56vfuo7P72ZlYQpDC1KKhZlZjoNerNWpq5Vv/X9fQdg9OFzuPe0++Wiaju4Ovv6HfwBOL6XMFiuJIiG3zLWbd1FtNnQTkqsreJvbWJq4w0a2SjWfZHZpg9GhXmZnorQ0OrhyYxzNbmNxZhqbv5XNyCyNrZ2ossSDO9dpaOvk63/wn1HcfgrJNdYzBmohwVZZpbnBt8dzNTI5ju5uxWuXmR6/jtrQQnhqlmBzE16vZ5ejlmA5ukZXdzvRpTDlSpWHEzN0d3ex8OgOBWHDKGWZmI3S1dbA9Ws3kFQbS3OT4G4iNX+Pu+EYDocdByVuP5zHJhtMzkbo6mx/smQrLMbHrmNIKktzU8juACvzC/ibQrhcnn3L4y+TaDRaPBSrIeHph8jOINWqQTkdJ5nf6wXlDwRoFC4aA54D73e57BRKFY6NjqBRYm55neEhLzaXh8jMHH5HmXOXP41DkcjFlvfcKyydVFnw5rkjSEKwHo+T3ojQ0DPKUG8z/V3NXLs1Q8ebZx/fwczEQ+z+LqqGRXx1lerpkf1CATWfETvFis7oyBB2RcIbbGN0eJBC0oa+ajE40E92c5OKUSGeN3jzjSNIkuDt775NYr1CqO8oQ73NdDUqjC8/mXpLkkQwGMTd2IHPY+fa7Cw9/aOAxupCmIHjrfQPHWNwoIHE1jpHjh3FLRuM3bwPoRa6+48wNDiI0dHE2P0FZD3L+Tc+jU0G484Nknkdt6+Z46PDzzze0R/q4PjoMAida7cesDQXo+/4Wboaau+m9HIEgI1Mgbc+daHWvrGtnfs3ogv0HjtNX7OPJpfO/DO88xuauzl2ZAisCtfuTDLQFqDR00bQ7z74hm1sDjfBQAOdHW0HT7EliZbmJlbXtyjn8uiWwOYIcOL4KKokkfrud4htRvB1jjA80Iro7+Dtq49od0scGT1Gd5Obu1e+gd3XRVW3SG9sUDYEru0jOM3iFpFYnqOBKg6bRCQaJxAI0tnZwf4dNy+fQ6EsLCHT3dtDyGWjp7cXh11jAWCXZ/+O87VlIUnSrgEsMXLyAuVClvGr36Hn2Bl8gRA9PT0ADA5r3B27suM0Je87kFbs3T8gS9vXtq9K0j53aiHZ6OntwaNK9PT2ocnmtiRP0pq6jgCOnb1MMZdi7Pvf4eiFN1E0bdufWcb2dO889UxaloW8vRYvSdLTP+/B4fTu1Lmvf4jq+iyqVnNIUxRl+636xP94Jy/pqf9u10MIsDkc+32vd6E+rovYJe++p/Kp9pWeJLAsgSLLO9efSCdA1Jyd9pTzLg6Pj+WGJ/c+zuuge/ObEe5Gcpw5NkB8fVuJ7ZKvdo94Mta2x4KkqE+c/bbHgnd7LDh3uaILy6KxuX27X3qwaXbGr8aeKc/L5tWZ57wDfcNHmJ+YIJ5IsrkV2xXnodbzNpeH5OYSiVSGqbu3SBV3GTuFRWRxnlgqi8Nuw5KdBB0QWdkgEd8iWyjT2dbEgwdTLEcjRFdiewuXNTw2i9mFCAtzk6SyBoHWPuJLk0SiUe7cukPv6O6Zg8TQ8CBTjyZJJJNsxp8Y5TzBRmKRWZaXl3gwMQvCZHF+jmSmgFNTD/ym3clVsdPglJmYnWd++hE2fxOhtl42FydZXlnh4cQCylMHKDu9blaji2RyRbpbG5laiJJMxElmnrWB7onSWwrPEF1Z4cG9B3T0DdDT1szd+xMshRfYLEk0et77rsiewWGm790hGl1mdTO+014NHjtTc4uEF2aIp5/YGVq7elmcfMDKygoT02EUWaLJ52BqZp7I4iyRlfiB5WheH7HVBZLp7J7rDU2NLE5PEI0sMrtQiz1hU6osrawdGEpAWLWt+8nYOhuJDACWnmZiao5oeI6yzUdTSy+p6BThpSh3bozRc3R0Tx6DI0NMPZyojYVYfI/xUvW0oFUTrG3GiG1uUqwaeN0wv7S8Z9v7q8Kh8eCsloskUxnsbi8Br5tSsYTTaadUMXA5NbKpJKZsIzI/x8mzZ59shBKCQj5DNl/C5fHj97oQwiKVSFA1BQ2NjWiKTC6Toli1CPg8qJp9z4MnLJNkIgE2B26HhsPhwKiWSSTTuH0BPC7HU9IKysU8qUwetzeA12WnVK7icjko5bNk8iV8fh+KoqKX8uSKZdy+AD6Xg2KxhNPtQhhVyga4HBqlYgG7042ERTqZwMBGqMGPJEnolRKJVAZfIIgiSdjtT77Ra/WMozq9+NwOcukU+bJOIBhEkyx0bDg0ZTt/FxJQKpWgEGdqw6Cr2YXd7cPvcQGCfCZNoWLQ2NiIKks7su5RUULUrructT5yu2rXSmXcLue2vGlcHj+aDDaHE1kSpBMJTNmGx+XAbtcolSq4XE4qpQKpTA5/IIgsy2g2hVQigYmC2+XA4XRS3inHoliq4HY5SCcToDoI+Dy7RBPkMilKVQuv24nd5ULoFeLJDKGmpic2gl11yKYTVE0Fj8eJ3W5Hr1TQqyUKZZNQqBFFljD0ColECpfXj9ftpFoqIWmO7b0dgnKxQDqTw+nx4/M493y2CcsgHk8gJJWGxiCKMNmKJfA3hHBor87E/2Pn7i22/extB+zKrPP8FGNRpmMSZ492vWxR6rwifOzcvSVJqiuKDwFnqJPTje+ers4ni4+Vsqjz4SBJ8jvZLet8QjkUBs46deq8fA6dssgl1tlMHxC5WVgsLix99AK9KIQgvBBBCEE6nXkRBZBO7YqYLgxSmZpnqP4uwXDeMVfLJPPM1Zb3h6XnCK9svXvCPYIIMun0gW7nRqW4E8T3hSKsF9R3L4dDoywsy0TXdQqZJOlCBSEEpmGg68a2+6/FxtomUFu/1nUd07K277WwTHMnbe3/9R234f1lWZi70hiGjmGYCCF2lfv4frEtW5VqtYppWdv370qzq0zrWXHgD0izsbaBwCKdyu6rl7X973EdauH3xE4aw3y3B17w6P6uaFVWiftTYfRimkdTi9v1PUhMUZPBtBA7bVWra82V3iSdziFETb4ded+lzR+3805/7qqLqZfYiB3w0AmBZVm7+sfabr9av6dTGQRP0jzO2ygXyRV1xK5+th73q2EcKKOwrB2XdbFd7p622L5m7cqvppCz+/r2cVrTMPbI/Xi8vqocCpuFUUrzvWvj+AN+EmtRes62sRGZZn49g10RYA9y4dQgAJZe4saNm2hOD/lcjpMXX2dz6hbrRYlgQ4jhTj/jj+ZxOWzosptLZ4/t876xd48AABpASURBVH8J37vBQk6iwSUTiyVpaGqiWsjSf+ISrV64d38KIarInjZOD7dx/fpNvD4P9x/O8IUf/CFmbn4fxR9CU8BQPFw6M8rc9EOKVYtUweCzb1zYH6UJi5nJh5R1k3RJ8JnXn8RLWFtZp7u7hbGrV1FdPvRyGsPRTouaIzB4lhaPyuTta3SffZPC2iLriRypeIILn/4BfNp7eR8IEhtrhBeX8fk99He3PfWz4P6taxiKk3w2x5nLr/Pw7W8heRuxq1CVXFw6NcT62hZNLoOvX5+kp6OJeDyGx+tHUwSKp4Wzxwb2lVzdVlKWUcQR6udYbyPXrlzD7vFTLSbB23ugvN/6o6/Q0NlDOZekIjkIel2k81U++6nLrK2s09Xbxdf/8A9o7OkDo4w71EOvs0Ss2oi1PsHdTZ02n41YPEGgsQmrkqd14CT97Q17Sqpk1ni4anDheC+p1Xk2dB9mMkwFjUIuy/Fzl5m/9X10hw+nJlMybbx+8SRrK+v09LQxPfGQimGRKcOnXzvDt7/6R/jau9DzSYrCQYPPRSZX4q233njlwuk95lDMLMIzU4xeeIPz584xOtCBQDAX3eTN1y5z8dJlpEKc4vbur/jKAsGeY5w/f47XLx5nenIOs2oxevIMZ44PMfPoIS1dfbR3dJFaW8E88O0pc+zEac5fuITqtHPxwnkunR5hfT2GbHMxMjxAZ1cv2a0N9GIMxdfBiZNnGB7sJej3IMlOLly6yPkLlzAraQQSvf1DtLe1Q6nAQZtaJUmmb2CQ9vYOjEJu387DYiKK2tjPhfPnuHByeOct9zTN7d10d3TQ3aCxFis9s00Pvl0i1NJGV1cvAz1t+4ycZnGd1Qx0tLfR2WBnLryFJDl26iobWaxdknd2D3Pu3DlaA06GTl3kwqXLVFKbB8qjufwMDfbR1dNPam2VzGYEX9dRLpw/x/kTg888cMnpbuTcubNcOHcUu7eFc+fO0WgXVHZ1rMvXxMXz57h46QKZ5JPyhZAZPnKCcxcuojrsXLp4novnThLf2C+jI9CBnllDCEFkNU53o8RyskpHexvdLX7mFlYxLRsXLl/i3PmLOKQS+vYMUZIV+geHan2br/Wt5gxw7txZLl86heIMcu7cWdp9GvkPaff0i+BQKItq1cSh1bzlVU1DouZ1WxvMEqos70zdDcNA2/aTllU7wtCRbHbs20uqumGiKrWp5KnzZw/0wZcUFVWt5WG3Py6vFiV6cWKcxbU4pmVhGhaap43y1hz3HzygoaUbVQLV4XziFCZJFJOrjN2domqYmM/YTZjdinL74Ry6YWIZ1j5lYVSraPZaDE3Fpu2LTm2aJpZe4vrVG+TLFUzTeqZC2RYLIe3yhTWNA1zd92JVy8g2O0IIXE3dHOlrQtmOGVrLVN7tBIptO+anoti2I27vCme9GyGYunuLla3UdruaGNUqdq3mYKZo9mcOVJvDse3eL6NtOzHt8jAHQHM6twfL3jaTZBnbdhna436WJBAH9JEk0Rm0s7QRQ1c82KkiqzaEENj9LRwb6kCxO3YdFyDtyJBaCzP+aB7dNDG3dx3bHI5aH0oyds0GSLXme569/S+JQ6Esuns7eXh/gnwuy9xsGJAIue1MR9ZIbK6Q0iVc28ok1NHD0swj0pksj+6O097ftysnid7ebja20vh8PhRFes9LhOlUjlBTE6JaoPjYEChq+wOEMA+MRVAt5LC5ArjtMqlc/oAUUM7nsLsDODVI5fYbcD2hTuJLM2RzeWYmZzCFwO9zsxyJkkluMTO7hDB1KoZEg99LMl2LnxFbWSKVPyj8uITHbjG1uEwum+H2zXv0D/QhqyqFfIrSrq3gj1H9XWjVJDanG4dNQXoX5fJeyGYLhJpCVAtpSib4mztZXZgim88zNTH7SizldgyOcP/Kd2jr7Uf1tmI38yh2F067jQM2vexQymdxeII4VUg/48jF3YzduPlKHnF4aDw4c6kYq1sp2tvasNkdODSVzdUl8lWJnp4ubLJEKpUh2BCgUswSia7R2NpJKOAhl05j9/rQFBkQZBIx1raSNLa00dzg31dWMZtBcXmxqzLJVJKGYAOWUSZbtPC5VcKLYVyBZtx2hdTqAmV3G10hH/HIBCmth+4GG4GGIBKQSqUIBAJsri5RMFSaGnx4vN59MwMhLNaXlygLjVDQi9frJZ1KEwgGSD9Vr1CTh+lwjtfPjbC5tky2ZNHcGMATCFBMxViLZejubMWSnYhKFsXpw2Xfb54SQrC5GiWVL9Pe1YPf7QAEyc01MhWJ3q62fbYVUy8TiSyB6qKnu4NcJvOkrukUfp+PTKaAz2WjoEv4PA5ymRR2bwBNhlQyTbAhuE8Wo1oiHF4i0NyBXRH4fD5K+QzRlXWa27uwyeDxPLWLVAhSqQyBhgDCKJMtWQS8LrLpFG5fgGz6SfsFGgIgLFKZHD6HStGyoZklLLsHl6bs9LMwdTL5MoFdBwLtLi+2FaOxuRlZAsusEglHsGQ73d1dFLMZ/NttkUmn8PgDZFMZAkEfa8sRKjgIBTzbfbstk1klna8S9HvIZ9NoLhf3xh9y8eKHG+Pzg/Kxc/d+GUSnx9nUXbT4ncTWlmkbPkt7w4sNDyKqSa492OSN86PvnrjOoUIIg3LZwul8Oi7Ly+Vj5+79MugaOUMwk6JUNRk9fXHfMYEvBJufM8ffOVZDncOJJKk4Dz518aVTVxYfEEmS8AYaOGDS+gLLVHA5XsXwKHU+zhwKA2edOnVePh8fZbEryOuLwjQPXu14J1Kbq+Q/ggjbQliUSrUVDPMZQXR2/2bqFSofwK374AIsVlfWMaslNjZfbDTzx1TzKbZS+1cYLFNnbe29uYiXSqXnikp+ELUgw/v9Woxqmep7CL77fsbYR8XHR1lgsrK8vvPXh71eLYTF1NTMe74vsRYlV/1wlcXB7sgGq2tbmOUUs+GDHZ+EUWZ6LgJAJZsg/l5OdD4ovwOuLIWXMStFVtYPjmL1rnm+x37Ts0nWE/uXmoVRJbq09p7yWlte3anTe5VDwtoz/h5TSG6RLjx/1KvZqelnOqC9bA6FzcKqFrhy9SYOj4dsfJPe02+QWJ7n4sULIAR374xx8uwFUskU2biNe1NLOOwqzZ0D9LYfsNAjLP7sq3+Mp7kVYVRp6BhiqNPPjes3Ue1OShWTS5cvMXv/BmVLBdlGX1crkw8mMCUboz0hvnPlFv6Aj4HhYcKRDS6ePYpVjjM+m+JEfwPXbj3E7XaxEY1yYfjCgfUqpjcZn1hAU8AZbKfNrbOlezjS6WdsfIZLF45z99YtLNlGuQqvvX6OsW//ObLLS3NnH24rzfxqCk1VGDl2lHQyw2p5k6mFNHa7TGfIwf2HM1hmBW/LIA1yhqlHs6g2jXZbnqzioyEb49a9KRx2DV1y8vqFE3z/G19HCzQiCwNXYxcnhg84WE8I7ty+w5lz51Bkibu3b3Ds7N56CrPM3fGHmMJEdoc4d7SPb/7xVwm0tVPM5bA5HGg2lYrQeOPiKZbnJlhJFLApKsdOnWRqfAxD1igVSpx97Q18jmcPV6OS4+79KYRZxd3cx5HOAJvLC9xSdUr5LH3HL9DsMhi78wiHXaOCgzcvnmLs+99BaE4a23rIJtL09le4fuMGit2JzRXg9LHh/eEwheDRraskqjJOTcGQnLx2/hipZJpydosbd2dwOTWCrd0EqhkKSvOBMiej08S1DoZbvWxGJsnJAaYfTVAyTYaHj+JxvlqP56slzTOITD+k9/RluoMOIg9vULIEul5zi5Wk2incIDB0g0ohj9PfzOmj/ajKs42Ass3DxYsXkawq124/wFFYpmX4DAMtXtJrC0wvrlHIlxg+fZFGvwdZEnR2dHHy2BB6LoHmDHLp0nksPces/thFV2CYJrOTE5y4/CYhp8K9cvIZ00rBxMQkoycv4bZJXL86xrEf+BTLY9e5smxw6uIbpFbnkHwdnOhrYXlqnKWtEpWKxac+ewkFk7evzPHWW28gSRKWXsYwTFrbOuixmujvakEIwekzpzFNnTu3Jxg5P0pXl87IQCfZyCNMSTA9OcWJi28QdMgs3LvOclpHoHHh4kUUSXDtxg046BROSUI3nrwxDWP/21OS7Zw8cxrDMLhz6x6CPlS7lwvnL5BYmSRc9HN+pIPbV66i6yUiWwXeev0ikiSRXp9DCfZydqQTs5Tgxr0p3rx84pn9qWiePXWlM4AnEOL8+Qsgqnzv+7dIOU2OX3idBqdC+P51llIVykWd19/8LJoicWN5CWHpVHSZ8+dO4XZoB8fNlSSqJYOTF94g6FQZv3WNogmGbqCXC6iuIKdOH0FTVWKzG5jP2jxnmjtnjwjLBM1Be3snp06drEf3fr8UywYdzppLrN3loszeuN5i1269pu4RlK1V7t0ew9vax5Hetv0ZAg63p+ZwtO0GXCpXCbo0QMLhdKFvlXjtzbeYn51heiLPuQt735pen39/CHzLwhJQqVq47Qog4XS7nxmouVjIsRoNowDtPX2ARCjgYnExhceusFHMk0rmWbDyYA/S7bOx5Q3U4oMaJrKiPDMMP0KwNPOAeAmcmkKhdPBUWDcsnJoMSPjcThKFKna3p1aG4B2jd+8qbE8fPGYzOkd4K4/XZSedrX3PO1xuJAlkWcXpsCEBsiSwjCqKzb5TH71cwulqRKKmCKg+e58LwPLcIzbzJi67Sr5Y237udHm2xVeR0anq4NzuF5/bxUahit3jR921cUvWPLx26RSzM4/IGzYunzt5YBPIdid2VYFtV/PHny3epl5OKJs8vHsbR7Cdg+cUB7Sg9eraKh5zKGwWHR3NzMyGqVTKtRgPgEs2iGXyZJNbLK8+iaBdKOTQvI2MHh1ha2X52Zk+RWd3B7NTs5TLJWbmFmntCJHOFOgZGCJoM0nlqxhGiUq1FsL/8QiSFDt6oeYevTg3j25YtDYHmFtcpVIushRZecYgkOhob0d1BhgcHKS1pYFqPsFKXuHz5wa4O7FAQ2s3CtA3MEh3ZzvO3V6Yig3VKrMWz1Aq5Hc2Lck2lVIhh26abGwkGRwepjnopmoKJFmhUinszMoA2pqDTM9FKZUKTEUTdLY8v0OZRxFspfPkUnGWV2P7ft9Y26Krb5COloadk9ieFeNetnuwikni6RzFQh53UyfrkTmKpTLh6QcEu3rfUZaNtQQDw8M0N3iobm8i21gNky2UiK3MYw900NEeYmpmiVKpwEQ0Tnfrfl8VU69QrMLQkVEq6TgHmoDfwZ5RKuaRHT5GR0dIrK++owJw+bwk1tcol4rMz4YBsMkG2WLlldyufihOJHN6G7AZOaKrm3g8TmRXkNHBHlbCi+QrgsGhfrxeL5qmYVcF4XCETK7CsRPHsKkH60ObZsPjrUV+1mx2Gpra8Gom4aUVmjoH6GjyE1tfZmVtE39rD53NAXwejcjyBqHmZux2B26XAySFoNdOeGkZb1MHraEGWju7MXIxVjcSDI4cxef1HLjtOBhqoZqNsby2gerwgKnT1dOL2xdANkr4Qm2EPDbC4SWKVUFDMIDDbsPtrc2KWtva2FqNspnM0BBqwuW04w02IulZUnmd4aEeIguLSI4Afd3NuD0+NLnKZjJPKBTC4XLR0tqGKKZYWY8xePQkfqeGpmm4H7eNpuHxHHx4U6i5ibWlRbIlk4GhAXxeD3ZNw+P1otkd9PR1sh4NU7ZsDA1243a5a/l53UiKgsNR21dh0zTcHh8d7S2sRiMk0nma2jpp8mmEI0s4gh0MdTcfOIuSZAW700lPTyuRxUXQfPR3t+Bye2hqbiS2vkZZcnH8SB/eYBNSOcXyWoyB0RMEtuvq8XqQoCaH28HyUpitWJK+kaN4Xfb9FZckVJuG2+NGliVsNg23x4PDruHQZMLhMKlMkdHjx3A6HDhcbhy2/eNQdfqw6VmW12N09A3SEPDT3tFEeH4Rpzf4SkX3jkajxUPn7r0ZniCttTHS0fDuievUqfOhcCjdvYOtvXjlV8tvvk6dTwKHTlloTjd1VVGnzkfPoTBw1qlT5+VzOJWFEMRjiZ3Ap897z7PcoD+OCCGIxd+fF+XLQAjxyi8dftI5nMoCi9npBcxKfueA23fHZHpy7oVK9aoxOzf7skV4LoQQzM3O15XFK86hsFkIs8z4+AMsYeFu7ORo/7ajlQDTsBBmhds3byNUDb1cpH3oJLmtZY6dOIEiSUw8vMvwsZO1cPCFDFdujOP2utErFUbPXKTBY98up8r47TtYkozmaeRIl5/J5RynR3t4eP8hR06c3Im2tbWySHgtganrHDl9AaeV49HUIqZRoX3wJN3NvsfSE5mdYCNVRHO6OTE6yL07txGyiiU7OHfmJFN3b1IVMnq1gs3pwjJNqlWL85cusjJ1j3jJAFNHsdkRlkmlXOXM5dfQjDzj9x8hywqKq4Gzx4dYj8wQ3khjU2SyZRNhGTy6N07JAN2UOHf+3M4ynqmXuDt+DyGrNLZ102jXeTS3jCIJGtr6GOoO8b0/+zauQBC9UmHwxDlEZpXwehIZweDxM9jKcSbmV8Ay6Bk+QYtP4ebNcRS7nVI2w8jFt9hYnOXUqZNIwP0Hdzl54iTTjx5QqBgIm4eTA23cuzNOoWJw7OgImiojLJ3pqUnKVZOllRg/9ENfQH0FQut9kjkUykKS7Zw9fwGwuHHtNmJbWQjLpFgss744ha97lJGOIEuPbpCrGhQKhW0PRCgW8gigkC8iLANLdnLhwkWsapartx7yqTfPA7A0eZfGwdP0Nji4ff0q+kAfruoit2/HCbb1Y9s+ZVuYVaYjW7z5xmXMcpobdyd487XTnL/QAFaFG2MTdDfXwqJZlSRLcYNPvX4RCYg8uknjwCn6m9ysLzxifjVBNp7mzOf/Ak6rwJ9+7x4/+Pk32Zy/z/JWnmIqTd/p12h2y/zpt77LX/rCX6C0McNcNIWcnGLgxCWaPDamb19lLd3O/EqCt958HcnS+dNvfZvE6jymp50Lw53kY0s8nI5w4UQ/AIsT92gdPk1n0AkIvv+97/L6W5+puXm//TY9HQ1UdYVPX7iIVUkwNhHBoyfoHj5NR4MXELw9Psdrb34a2apw5do98h6TrhMX6fRr3H/7m1QMQT7/ZKNXoZBHQubI8dMA3Lx2A8V1hK6OLk6dHN2Z6kqyjdFjp1hbmMB+/FRdUbwCHAplkdyIML20hd2mEE/t32GYy5VoaHMDEm5/gMKe+azYt4PQ6wvUXI41N5L1ZHtzMp2mXJkkEQHsPmyKRHdvN7//J2/z106f3/E9tIwKydg6d8fHAWjv7GBp9iGbmQqqLCiUn5Rn5JI4fA0792ZzZXpHXIBEwO9ndb2A6vLhUGUkU8HnqzlcqTYF0zCRHW5cdhtIFl6/D1mSsGk2zIxBtWLic9Xc4EMBD5uJDDabHVmSELKK1+ehmMvjb2xHApzeIMZ8eEe2TK5Cp9+x87csydvRqSVcqg3dEHgDwVpbqRrCMjl+4TILs1O8PZHj2JlzZOLr3L9ba4emtjayG2G6vDW3eW8g8JSrdK0vKoUkt+5N43Q6iK4lOHvgB4igWkwTjld57WLLAb/X+ag5FDaLpcUVRk+c5uhI/4EGzVBTkOjKBqZpsL68jAU4sMiVq1RKedbX9hr61lejVA2DbGwZ1fNkIHZ1tmP3tnDq9GlOHB9Bky3uPpznh//Sp7l3f2JH6cg2F8FgAyNHT3Dq5Em620OsrCY5feYMA13NO+7GALZAO9nNCBW9dmpXR0cTswsrGIZBJLpKc1vDszyg35VQg4fIahzD0JlfTdDRGcKo5ClVdSqFNPFElsaWVtaWo+iGwXp0EV9r6879bS1+5sIbGIaBbphoiiCZL1MtF0hXDewHeB3quknf0FFO9IcIL23R2NRC38hRTp06xUBvOy1NXiKrCUzDYHW55upuswyKFZ1yPsXmZpr02jLBziOcPH4UVdo+W4OaDI/bWAiL+/cnOHHyeO10srpB46VzKNy9Gxr9zE7PkC2Z9Pa04/d5QYA/4AVZpbWji2p6g6WVdSRVRXUFOTLQzszUNIlUjvbubhoagkgCPC4b8VSefDZFugSnT4zsRNp2B5rR02tEoivkygYuxcDV1E1TQxDVKKK4fNgUGUmSaQn5mZudY3Mrht3jp6XRzczcAobiobu9Aa+3FmhPkjVCPo2ZuQWS2SLd/SOYmXXC0VXcjZ30tjWCEPgC/u2TJmQCfi9CgM3hxqmpeHy+7Y1dtdmIQCCpTrq7ukitR1heXaetf5TmgJdQwMPs7DypfJXB/j5CzW1oVoH58BLC0cCR/vYdt2lvQwvF+DKR6Cqm4mBkoJeF2Sk2YimOHDuB225DAP5Azf4ikClltliIRMlWZI4e6aervZWFuRnWN7eQNBcdXT2k18KsrG8hSeBt7qSvLcDM9AzJXIWu7k46e3vZis6zmczS3dtDMOjH61KZmY8SaAxhU2TMSpHV9Ri5bIqtWJpQSxNy/VPkpXEo3b3fjcTqLFtmkNHupgN/r+YSPFhIcv700Ecs2SePyKPbyJ3H6A68ohFo6zw3h9Ld+93wBFtRxbN9PFWHh95u20co0SeXUGcvkqve1h8XPnbKwu7yccA+wR1km51QwzulqPNh4Ql8bCasdTgkBs46deq8fOrKok6dOs9FXVnUqVPnuagrizp16jwXdWVRp06d56KuLOrUqfNc1JVFnTr/fzt1bMMgDABAUESRqJg3MzCb2caVqbLCd1DcTfDVk5gFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkJgFkHzWWvPpCODd7vue3+u6zm3bfvu+H08HAe+z1ppjjPMPOMBgs3W0FK0AAAAASUVORK5CYII="}]}