{"current-slide":0, "aspect-ratio":-1, "slides": [{"background-color":"linear-gradient(to bottom, #d1ff82 0%, #3a9104 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/diamond-upholstery.png" , "items": [ {"x": -547,"y": 721,"w": 2521,"h": 472,"type":"text","text": "","text-data": "%s","font": "open sans","color": "#ffffff","font-size": 42, "font-style":"regular", "justification": 0 }, {"x": -535,"y": 1085,"w": 2394,"h": 315,"type":"text","text": "","text-data": "%s","font": "open sans","color": "#ffffff","font-size": 28, "font-style":"regular", "justification": 0 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nMS9y5IkybKu9au5R1ZVX9a+MQA5MxABEWBwXgARxkx4Ah7jCA/ABIRXZMAI4ey11+quqsyMzAg3Uwaqv6qah0dmVq91hGyprsq4uJt9pqamNzOX//C//S//03/z3/1X/+ef/vTLv1MdkAY0adLHUKgAbQBQQIEmqyi6QhuGdm2tCQBAgNEV/BGI/b/BvgtAFRABdCikCRQDggWCJoqB0ftoq8r55bl//vzTopsoBJAmImhQHRA0+57YbcdQtCYQEfRtqAhEmmCMoa0tAlUoAFWFaENb7Yujd1WoNlm8qQOtNRmbKlvst8BVn1SaYNWfBSqiGCoCNFmkj26MZAACZ7TcYaQY3Rmo3XZipAKF2mWUjBQCgWARxdAxurZV5Xx+7p8//7zoBmfURCD2PcjEiLx/jJFi9BGMpAGKPSONe1z1cSytSTNGfv89ow4Rgb7FCIoxdoxEfCx2jOL+6hJn1xxjaFtVns/P/cunnxft9gW7xy0jVZNtWQRQweg7RtJ4d8CIYH0Q0a4YY2IkiqGtNembql07x+Gi38faVmn609uMmkBHMlJt0DuMoC5F0gDRA0ZIdjeMhpzPL/3zp5/eZfT47fz//N//1//7H9b/8r/+z//3f/8//st/i+snu6E3IP4tdiMEMZ8cQHmfDc/BsxGon/HXFfN9qG1aB5YrMP7Brq8N6Ke8r+jue/xb87b80Ta3q3V/bQBjMQVYP18vEP0ewOkVwKds9/XzLaPaZy3X+wij6XXN61VG0bTCqP+j/Xss9qe2R9T6GuOAcp//PxjFDd9hNPz9DzAiFxwx2oBlO2bE70i5XjDi/feMSrv+MKMXAP9ZXudmrv0RRvUzu/FtCoyPMPonZ7QCoxWZ0Lw2FNB//geo/B/rz//w07+DdOjpDFy+pMBFh4vgseE3jecgjDIIyNfHvhG767UtrxmwuQxzUFoqkYDT/O8y6GxHXIf/9IGVbYaszd+TvIYMYH11UEhBOZ2B6xfkxC6D8Saj0rfKKISicq6M2J/KCDM3FQCVDftZGKW99EFGvfTniJF/f33JNpHR+gJsn8s9/Dt1Ut0w2snLxKgsNpVR7eMRI/alXX3ilL4IJ32ZnHUMY3Eaeb+/mZH3pW3ACmD7NDOaFECVr9q2yqjI3TQXGzDeYLRci0yQ0QUYn3zO3TISKH769fO/a6oDOsS++PCcNxni2oYtHv672HvsxMi2YDT7ww7UCUKlUTs/HDAFfHDg/FrLNQeb96/XVh8ENkD9XrLtPrebtMNf4/0B/96w309nH1/N99iG0xEjDuZIZlNfyqAeMsIdRoDeMGo7Rhfr70cY6UcZ4R1GahxU8tpkJB1Yz6W/hTdKHydGOrc7GFV+yAm6Y5RtJKOlfHcxxS/9DiPkHzKizPJ+e0Z1XO8xkhGMbuRINlcihZFWRrhlhPcYtZkRFUKVI+kpAzeMXmY517wXVeLa2iJaV8f1DFx/sptHvKJqdwqed66NYjlULan5Xf7IQFoBao1vG9DX2/e0AX2x1UokO49ipXA15WQUQvZVDmWQOmGyMQdmJ9QUxfD3xwJtowjJe4wyvgMiHi3N4ckd268W9xmp7BkV4dHFLQw4I1/ZOPGl22dGWcH/LoxcqDotv8KIK+r1yx1G7QOM6mf4V7XOCqO2uTIgI/adjNZ3GI2/E6PSpvVlYjTJ0WhuYQyz5tUZVddlz/1NRvXzlKvu3MjoCoW+wWixhVlPRXElI5WBdehmlgVNMvHJsH0G1MJrygvWOAYHixOLr4dpJ7CAZJnUQdkHIVbEnpqRioID2RdfBRdgnGYLIQbIFUUopqKFRV0IRlE4XKlsYosMe3l9LZOY3/H2xyBxMvwII2pr/65IYSRvMNqKkqqMvK/S7XPdFcZYEOZwMKrBryrle0btgFGupD/EqCqM7dPbjCblWRnV16uSYPv99WXL7x0yKnLUNpss/8kYqY3l+rJj1P2fhRGvtb4A/VNO0ENGuCNHWvjsGRVOy1b69h6jqy1MSEaiAh2ClV/U6LyvAusZsn2ChqlWLAlFTLRy1xxIXz0UIycxYQE+CTS1/M4q0cZGwgfWTahl+GCXVbncPmG1bF8sxPU7pa3s++kM1aVerAgGrR3X5oC1Nxg1hE86MUJq8Lhvy2uTUbQPMUDGqHCvjCBQISO/L83MpsigZ12VSxtCMdX39WOMxoIInFkDso1hTTZv5wYsA9KPGHXvl/c52njLCPcYLSXWNTGyvqlPNKH8jmYLTxs7RnNfQzncMHyHEQCsZFSg13Gc+ugLAhTSH1zWDhjVPh8xmpQf5s9XRmF1vMOobSa3zkgBiIisKgMqpm1UBiR8H4Uubkqqdz58GuTgxN8UPrHPV7egBnH2waopus3OIxoJ2RwiXZKeCiSUboHHe09w6ufK63zrdM4VBBT05s20AbP5sWc0nNFPzsiVYzDCBxhpfncy/Sqj/FoIgit3M156YUQl8wFG+AAj9uOhMNLKqM+MQo4EwOKMXosckVHxtyujcGnvMBrNm01XhDGdVhhRxqoc7Rm5RVFX4TpGtR1vMkLKW5WjagGp3mHUYry1XdxSPWBU73nEKOZUZTRc2RRG+KOMAGmCtUnz4MfIL7GzYW5bBkBGu1mkrB80gbj6Sr6tZRVrHWGKAYhVuCqUGhkXXyXZCbosfk9VuBkPQJlbFlfk1RzLNpnRr/Z9moE06bUBcOUkm8HtLvC0uiZGvprTJTlihKK1d4y0CBO0+Rzfst83jPABRgxkkZGkqDujGJ+PMMJI//tdRu0+o8XN7Y8wQmXESVEYMaMVKVHJFVbZv6pkjxhtgK7mKh8y8mZM7qG1hdId9QjMnk2MRvYdzcdzL0dl4bzLKBXVxEhzodUoYiIjhbarfVYLo2CZMhAW+CEji2GIK5lVhwHS0KbFjB+uqZYzZPuCMJmrRgVLQCRjAwU2CIf+91gLULa/l8sVc5L3H6vfR63h0u3SYzUzygEqBzhFMNvgUOwzptl1eSl9pjVQtHmsrEX4Rp28zqjZQMv2+ZYR2d5lxPcGRrtCRO8wmleCNxnpESNMjPLn78mouJ1ywKi9mkvyIUY+ye4yOqWy0toWTm7J3w8ZWSzMXM+lcDlixMsbI40J64zaS96jvHfD6EaJ7Rlt7nF/gBFjNFjiffsZGG1z42GZGUl+5qZ9HOOJ0QrIFaonjG3oarJSO7kgzVy/aNug6xly/ck7WwSEwgH1RlE7SfJuJU3n781uzN6HLqsd2+FCndq2e3kBg2rkqKlRKXA19iDDVqb1DPptszD0HIxogpqAsp+jMsqB1uUFstU6DHmfUby8+ZiX1SnMTrFYxORDHzDSYtFNjNaZUawwC1S6K+Ado3a1la4yCqXSixDzr8JIixzxA2QE/QFGIxiZh1AZbXcYvSNHwcjv3TbTce8xqnU+nBOVUbX2GGPbMbI+F87VkgJMsberjV7UqhRGKNc5YAQVKzcArY0do7jfXo7wBiPra1tVVmjzgAw1Wd81yAcaCj09msKY/DEKROl4VQbSPSZiKRvR5gHMEa6AaJqbYSNQiWAHlAILmNZrw1aJmmqLCQe7v7qzQrPtdMa0+tTUbywrvsKxRTT73mO0PkG2wogr7jTQhRHwBiN5gxFvXxR9BKuKor7HCCkYQ+hPp3Dq8vIBRtXn58rH94q1yL9pik+MOMHfZqRvMKKsBCMVy0zEgl7kaM9ImzNyi+xDjFzRrztG+hYjIKwCXrd2NxitUHTo+mxKtTKKfpTvT3JkyphjdctIi+z8CCPg/PrS19ZEgOGFI1V7VY2ck9UsjJ/ztaNUIVcfX8XFTRsL7Gjpp62gNsD0e3lvD2DFalU0e1gaK8wPLFqcHacf6GWv1jSFrs/2WkSTKRD8rs7aODIQGVR8k5HfY2LEzwgOGNkkOGak4TO/yQgzozCTyUgGFEXQtPRzYuTtX17+GKPI/OwstomRj8PijGIVP2IEZ7RBRc2KBG4Y4YhR3H6U699jdEK4bZM14JP9b2ZUXArKdCjfI0Zu3S0+16T2IS9VF5uw2v5ujOiOWXs+PXxa2gC/5JM99EIVdI0GQBW6PuZn1BtdK83QTTuiA+Pk8uyBIAUYiNIhnpql6erXCcW8QIcFoGLd8qCdNdU6rlColEpPtTZEx71oS5dz3DsBZfbFJuuS7wePslJ8iJGtnseMKKRkpDMjVEbyPqOxmGC8xWgsUIxkJIUR9wR4Bmdm1Hd9foNRmK+VW2G2Z4QBPT2/w8gWG7v8WubLAaOogpzl8ZbROGA0nFGfGeHvxQi7f4/S5yNGrkzQj+WI/auMFHnPO4ym6l/F24xUgZA9YPSuqylyQaZgvGGxEcVTLiFkrvXWZ8j2s8HaFUopsx4uPGZKK5gy4oqkAEQt16uinlUBACkLZongh4LgJXxyjQZtG7RdICzcipiFX299QvizKruVQPN1rmrRp1ZWCSACjcAbjDw19kOMfCXQY0ZDNMxIWibvMYq+B6MrtF3dPy+MNF2oQ0bx8wajeG89YESlXFZabWZRrWdzSdDtM1wxVdx/16KEcizIKOoEXA1IGXMUM3pmpDtGgKrxmBn5uB8xmqyfjzIig8pI3me0vED6F4RiCmtbLOU6xR3uM4IrymSE+4ygoXBsd4hgHUPjIqQnY0FG0CUjCeE/rWYaro9o20+RQgKGB6EEjKraTcVlzs3vElA1reamIeFRITj4sEh8MgSMalqP1dwa2SyKqwBN8LE+IVKRUB/4IlS8DqviIqDk9ZVcFQ4ZUVhvGals0OUJrX/5ACMgYyRlcnBsglEVyncYwaycZHSCiuXPRbkKLVAZ0PW8Y1TjCJVRnyb0m4zc6mOj94wkGD2j9c9gutYYXW2coiYEO0ZIRuJ7rLkYfYRRXFHKa3LASHeM9jGKes33GPEzbFup4H2T0RW66A2j0a4Zi3qLkZeKG6PFGRXDYFqENdo89QnAKjVtpAJWFaqvdrEy+SoU+tR9tb48om2/IIq7ogikx/c5IXISsqFi14lqPo33Nar3HGp5Xfze9hUNK0M8cq1yhejJgC7PXvzCNljbctYpLP2kxY9MpWW61jV8DD4VlZbfcxV6nxGFq/tgA8eM+HuDNr//xKgO+EcZUakOQE8AFGN5cl+3Mhp3GK3vMKJ5zgre+4wQjAb68oS2/eyMuJsWhVGxVqAzI90xqm2rVo6KG8/3GOmOkS+MGIUREJbkPUaai8B9RuLf+ggjizH05Qnt+gu0+X4hZS3GBxiNPaP8uWXkiqcwEhFZpSnf8xuwg2yI3zSyCwKlOeSR3r5+R+ue6on8rWQaMH6kXI+qtBdFpZg3wPA7bJYA6jEWoYlkb0bgxtOApo1fYTENDqZrSqnt5MXZlpbmd3xO814To8qt9lWg4FZ4U5hjfYT0T3mvYISdGXuPkZSVaZdpqN0Q53GXkefRpQN/N0aZSs5Co3cYqZiFFauYFkaVBQ4YtbjGISPZM8oFSsMaICN9h5G+zSiK5T7CiCUFJUPxUUber7E+QsZDmS+u8Lg/J34k73GXkcZt32VkbghykOk31Uhus0yDaNuZmuykreZ9eUbbfgHAoiANpSJeRVZNxEwFqv8O077uZwl2bkaM6ML5YNeGB5/EfCxWLY7To9+3CDyAeUWYJ67QjB0tT1EK4XCYEf1HDrbsGE0pLpigtQuwY2Qa/aOM1M16W3VEG6Ia8COMuBegBH7H6bvFeCYF5owis3HMiPUtxohtKIwimE1GI/sN2HfGntErsJzRtp+y/38zI/ahui73GHG1/0FG1dWjHOAeI35s+OJHRgiL7T6j1RkNtO2L34uMyLcy4twiI7tmMtr833tGezmydrVGC0IFsWtxiuRKaqNq5sQmk81AjgVjfQSgGF7bwAIWi8RX0x/2u8PNlA7cj/exqSY6tavKNG6WCRlTNmEsz5D+UDImbItfOKLC7hN7QEqLC7CPJkcbyCiu9wOMtE2MMDHylayYiIr7jELXvcUoFg7rDxmFe9Y/p1DtGWlhNG4Zmas633NiNPaMkIxqundiZJ8Zy3Nh1PDDjFAZyQEjz8bx92CkhVH/AUbrzEgro5SPtxnxTzLSiRGgco17jMXOXLnPqM6QGtAkI7X4zCEj4JaRYO06SnzFtJ/4mxnkpCbvcVEBYGkt1ggAGA2DJb2sm2cDImjnK81wrbUPSMWE9fsqLOjDQa0DF+3zDkvHaC8efBwBWNHQxkNabiWrE5pW2D+7roy6gkmB/yOM1O+vyUiAIa+QsWfElacnIw7gIaPSHoVbWDtG4dJQCKyKcrRXZ2T1A0OuwFuMWOBzl5GWMWMbMTMaKG7ae4wGhlx2jDib3mMkiJX+TUaKXHXuMNIGRbfUrFwhWCDj5Jfg9/9ejFjLQRdfQaVvjDZjUfp7K0eVUVFSdNvCAmE2pypeZ6TFwnJGXD7XpTWJSLsHeAb6DNb/L7BJKLqgtxfvaNHmXJWXM6R/Lo3lxLQOhZLgqs5BrigZXIkCGpp8Gp1X77+yUtSrDm3u0u+yiHtW4ElmFvwCGgEimuoHPqUP/i0jZizkgNFrCRLvGLUXyPj0LiOZGM2cfowRjFF7vc9oUs7eL1ccURQl9xiJKwQyIhVeS80XPpSjBRYLq4w6tJ2TUfG/k/URI04WTL9rpD/vMPK/bxhRYeqKIRsaFp/A7PeeEQPA2DHyCTswKf9kxOBo8/a4u4dWGOGA0UuJYRT58o1jfkS1zzXKz9TjmRGYKZRgxE+tQwdU0qRkB0PpTjlau+GQqytjrrDZCGpRbWe0/iUbdRP41FDMGdBZXDtTK1IkJJRCpOOkZxqIpqtPGPH8dN57MRMODRinFBgA3AAU2Q0HXn08+8nMzMxIwQDQMSMcMxJTGG18jgG+ZTR+gBHi9cpIKqP1iBH75XEVXdwVHDnnyEiOGMXyXa5Foa6MaDlpLOJDLn4dQMaekS8ADWihMOrqvGfEe+wYgSLsk/CAUaYT7zCK2oUFY2KkB4xoGbzFiD+V0ShyREayY5TyYUpTwVJ1Y9TimlQMEcycGJkCF800aiz8ikmZq4+d6CIrNWUMQJkkghbpREWLCat8T2lCyzRQcAU02hmt/5xgGGWN1Z2ZkPSXTGmZ36VYQlcNX0Xpf0c+XuERYp6i5YFRRVkVGoDVC6Fyc02mIhMyBzdWRLoZpe5kDhYxwErlCWhT8NEF7zKSF7TxU9x9ZrT8IKNeGHWwaE1VMdYnY4Q9IxQGq0XfBT/AaIlJo9BoS04PrvytfMYLxNSsDCrVW0a22g15Qes/Yy4aqnKkbzIClmjQESN8hBE+xkgxuwTJCDHB7zICLRIyusAm5wEjhb9ORq9o/Se3RtLqsTanEp8ZjcIIPh4NIwKfhdECtOEBP1WP2qpEL1QZGFPzbdsrGGDS1DCIwNAwzaRqg6gA+vLkrJniQWjcCAQpvOEeVFGYORcBJQHLgFVd43nfx/LswSy1FYKBoZE564Ds/jmDTtY3SwWz9BfRJpvkdj3cZ8T/nONor2A0ve63iQDjDSNFX578YpWRX90ZJKPlfUYYEF2TUTsbozrWdxm1H2SUgUEJRkhG3u6Z0TmvXzIJt4xgY0pG5bpTAFexY0Q5EshYC0NXLjeM1BktH2REOdKYrGSEu4zG+4xCvhp6O8cc+Rij4YxaYZQFX8eMZGJk80pK0JmMBNfXbTTzJOhzM4KLmOzxx33aAA/xWK/GzSOoSLjesN6e4pNg0MgjtDYnTPuG0kGuxuoTkiYS2wgA2/LdAfuAeIWjqnjpfAuhGj6Q0q1CT7FBufLHgPmfEPARk2EcMdIW7bPx2+wbwQgY/l8K1j1GzztG3CCH+K4xGu8z0h2j6JO6ZUhBOmLUgGDULc5AYcMRI437JyO+t2ufCka7xv1vGWHHCDE+Qzb05VwYLTFGvN+UEVCJ9ubfprwrI4ViWx4Lk48wWiyTIFdjNJYfZNSizYeM5OIXaj/MiIp4nmsfZKSFEa8Ls4Bfx7ex6oAyj2p1Dpw4NGHc3JXNAinSzUyJwI3fSEqBTQSHfDJKx7Y8Yuk/wY4/o8/l96CLwapNb30GsBih1fBPzaJgUHIUgPTrclDyfIgWnzFzVAE8QCeTrUaLD4JAwMyIAy8bLLd+2jEKRMi03z1GT87I2Xq25uOMalBSvXq1lAPvGNX235yhoW6OQgE9GSMdyADYW4yqHGncY8jFpGycUqYmRpqxmB0jqyfYCiO3smSLzxojBupKs9x0J6NwL2T8AUaUe+vXkOsbjDJ2cKu23mO0YojFjQSYWE9yvmM02hUqw+KFjDv8UUbe59FecFoe2tqaSBY/baEgKKwWGFQXJMXACJ9sKgcHshEucOaH5ZkMvZ2x9F+y4SEjNJckfo8AzuCuUp84cLO6fhYAU5hzcZentEZpJ00vLJaeE2Au3pK8rLJYB8g0aj9gVFeCPSOZ4auk0N1l9LMzon95wCgCYWTkCttHf7Rn0Bynn/+HGUELIwptZcTf7zNiKpKuB+Nertd2jJDKi9kOCERNyaQcYccIB4wy/jMzctfjhxgtfhsGl5v5+O2Cphz/yojXKynyCCpTKd5jpBMjaC1UJKRcQIJRd0bygmX87N/9AKPiMQQjKYwgWO05i75SScIQCAaurtFaBm0iiOM+IBSx+aSsolBLLxpyidVua25h+DVDk5fezM/tpAa0xveFQSifqAHdOj4igOnXYkxENpv4kQ7SED64uZkHzTQwcDe83FbuMrr4ve4xonWWjDi50hQudQHSsbUnLJ5JiiDpDSMgg2ncJo07jPR9RgAU9xhtfxsjubhbK7u+v8dICyON70E6enuMbFssWoeM4KNSah1koC/PP8CoBtc9Zc4FFArpD3aU3ThBpwl8xMiDrXwW7buMgKjFKIzEr6F3GW3o7cm3YewZpZVzywjJqCUjHeE8MeDIwEvDwJZCDPPV+BBZ8+EMXLg5Sr/MfG36eBE0QQpCb2eX7WGDUhoPKhaIC5H/G8DWLIBjWQCPKZQgbASIOHFMqad/p/QfvY1QwM00RQlY+cSxjvvWZNfIM6NrtG9mxODWjhFogvZgZJ9nnUBacN2tp/uMZMeofYAR7jNCZYQdI98dSpk4ZIRjRp5CZtOTUdsx0mTgCjAZIT5PRgpFby+hSG8Y6T1G4w4j/r1nxLEsjPi56UyS1YOe2+RuJqN2wMisc0uP3mOEIrNkxDG6ZSSF0UDHaPaclxGMKK8p61WejhnZfy1XQ2o627WpEcixslTxMmcKEicIShCQ/jUDJwxa0sRB0ZDb8g3MFqRZl3Xtdo+E0pfHyILECuAlvdM04mdQYiohbHMdPNusMSkv04SMCV5Nam+P+ZbDBPGGEXnsGPkqlYzY53uMvt9h1AojfZcRe8TPvs+IK/SOkcdijhnt3EIyUk1Gep9RTAhnpGQUf7T82ycwLBZ2y8j97h2jAVttmQWZGcmO0RoByxhHMhpkZPGZlH2zSIYvEPGZENA9o4Eur96WLP8+ZlSzKm5XUiEWRvV38UXfsiSphNNdylIEds8YPWemyO/VZMUq0qT6w9S2zPtSFOHmUZpjgJne1XtW1HyzAWSAiCZOGDPY2iPW8adotI+SD4qdF6E63Kxei1Lg9Wh+mxYN/27aMYvi61VTi34c/VorRBnoaLoGxNgUFGa5QFtHxmxyuh4xoskqKIMfjEa5P1dVjbapuyTr+NXaF4zGHUanGJmJUZ1MEH8vJ8ctI0UtyU6/lowGmiteVr/SnE5Gmw/n38Io2xxs/A8rblVMuJfxS2HEuFBlZJsdRT/KiKtsaIyJUciSx6TshwHFkf8GgHcZSZCgLCSjEdSyDWQExNzlWMLMDBVF8zjGkA3azljGz85ofJgRLY2uHWudQMMtCtHUnHQjhWYYAFa72Xe9VJou90hlAJTdlcGckXRTRlv7hqX/iizGAfIwj46tPaJxy3BcpNbem4AIDIxFeb0gCvTl6mYjE0uaayOiw1wZrhjYsOinmJzWF2tf99VSUBnJXUaceAL68UeMssqS/bPYgVVSbu27BfRY4ecxBfLvwWgcMAK4izHawKq9Eg+ZNxu9x+hi39bPSMNC/2ZG4BhCCyMqhzYx0sJIXU6W/nNhhCKj7r/rWiY7ZdEn4YcZ0YRHfA8YftgVA5pk1ND04ZDRJq+upGdG3IkaSitKx99j5H2QzMIMzgOPH2pjJqky4tWd0Vh3cQ273tJE1tZWgQq6vCIrySi0yAkT2pRaPVeKXIWpkdM8pX8GAE1XS1kWba0QtzB+SUl1zXddvqO5lkvtSgHg/Tq4Eoi6iT0dvrr7DnYrHYtv1AREPH/e8YrmCoPbsoe8Ilc1Xv+IkRWz3DLS8r3KqPvkMvN31JJh/1dvT7560kUwRtvyzQXyLUZsgwnkDSP9KCNTxjOjkzNyq6N9lNF9OYr+HTKy9s+MGMN49tWzWmzA1r4Ho2iTa6662t8yyjqImr1LRmVM1ZYlpnhlnFxhXF2Rw+VIMTzWImGRVEbZ7sqoWrfvM0JhREvFFElvZyzjJ1RrVqEzIypaancM9KG6jtHVFAUmUz8ivtEZTUVAcy122vWI5IJaSSU6RxEefkIVI77q/1IZuLZvOG3/CKZMt+Xb7Fvz6LTQwArVFsYZxdDHDaF0JLV2RJmRkXOzojZk2fHwCWsWhk0G8y0F4paMXT8HO4Xd2kIrQgujrB/QO4woiLeMTJFt7RvW7R92jNY3GAF82tbfzEg2sLS9MrJtAG6qygtEWygKfZNRmSATo5IZKYzy+z5JdoxoVW7tO9btT4XRdzOrCyNaZe8zovmQVpdotp1xEbiFEFsJsEB1oOnJ6h4YIxCXI13A/UK3jIAsaq+MrJ14h1Hy2DMCGMzf5BFr//XDjFSAJgvWgW5GSfjpitzFyHRgPe0K4Gpuuy9HCEcG5/i5DYwjRC0Gi09CO/J7Ddfld6zjV2ztu6/MdXWbrR0hsLIixoDGypj5/gtfhNgAACAASURBVNmvk1hxLVpdNXd3oVh963auhVkvT0ajMJpTUlyRkhGLaDJY9aOMFIrr8hXr+OWDjKqS/zFGLJZSbyMi7y/ZTl3R5epilTGpPaM8WKa6SWw3GWlh1KbPUplzEmi0nx69T19XWtflG9bxc2GU1gyYLaAi1p2COGKkG3hkXraJaV9+rycjLYzGii4XNM/61LGcGaWVlffg/1Neb+WIVkhh5POX6edjRt+xjC/o7fFDjIZ2tO+P364yVliq1HteDuWgdg3xn8wxdtzTc8IUWJoykyBTkCIFa5Fi2xptE+Zl/Y9g2XKmrzzGUWoDFEAc5e7XintoQRRSQIHle9mGOLlZ6UPbNWWs2OTs5wYs7zDS6GsEtohBxVJzEyO2jcHlI0ayY2TCcJ9RtikzMFJSmXY9OWREU9sYxSMiJkacwHtGz14ncMRoyXRkmQhxGlQwQqQTjxmNHaMx9SlTm6bwX9b/mLIQAfy3GGHq78yIcaI9o17aqMAUN9oxak+WSQpGJeCvS4zRLSO9w8gXqyNGZf9LMsKO0YbX9c+FEVIZ3TAyy6mtD63RNOJAAAmEvgsr+Ag3BgnqgiSmoer346bFdCtpI0Dj+ooNXZ6hClzlMe6d6auckAZsLsDJ/zpsJZRi8XgcRu3fLB6yNlDwqFUJH57/tj4PuXyQUYnIozDCO4xwxIh+uV9HNmzOaJOn2v1bFqFIajyCa/MRo5a8yQi6Y4SixOxrJjtkdH2DEXZyhANGrTAqE3OSIYn26k6ONBidoarY2nMCeouRzoxwyEgKI71lpP7ckbuM7P1kVCblISO6DmSAW0agEt8z4rX2MQ5TDCMYDWztPMlRxVQXGwFkXcQ7gWsJAikQ+2hr7ILD1eJzac7ahpMpDSQ9OmUxDgRgATMcNtgbz6Pwvl7bN5z6r9lo6W4aN/dx8zQst69Ad8bMsDLrA5YCNaINE64UBPU9I0vUUYivMsM/d8yoDNCOkQQjvcMog8rphnjcYc+oPce9VMjoT9GeY0Zb4UppICMgtzunGzUfXXfEaCuMFAhGV2d0epcR3mSkiKyJVkZACj7NbLosFkPb5DkntQxc5TtO41fz7/1YgLuMfPCU2aY/wIhyOeCM2mthtOSpZFxU3mSkhREmRuB5MPFE+3uMqgvYoaLoE6NuMYzxC8KFQWVk1936prZFXRd0XNCjdFnSNKOupZ/laRiaKVOlp3JlcoHWBu6Wq5aImbisghu4tkcPkHL7rWmzS3sMzWjbsV17Dlo4iHtqrDQaZmdaiGlVZF/4XbbLza2xoMsrBniqcjNDdKzO6HrACHcY2X3SND9iJIVRK9/p9xmBjAau8h6jcs9xwEgrI1upuDJyZTtm9BJ9nBjJazDSNxjhTUZ4hxHjFR3cdTxgLGIvEdjfjqs8heX4JiPcZ8Sx46S/x2i4dWGMzu4qtB2jF/TYUfweoxH36awyDgsQiCLsQ0YojOzfmzzdMBrYcJVn0GpnURhU7ImAUEgTWUVEoIKGT7FSNH3wZtfAl/lD5tdYBoGPAshpWaK6iukaNN/43AQqmE38vAsqFL8jO3uVR6z6s9kCCtAyYIoobuOaNH8ysq/xAYJnLYkpvWp6dbEDRyQCWvB+NzT9FBbHLSP6oJURg4dHjNjf+hppj4nRNVyOPSMLSm/yiEV/BvfUzIwoeEUpBCu9w6hhqrfhpPDvdbES4vwuwINT2njwSliNAGwwko8wquN4j9EojGzSbe0RXEGhKP32Ogx5wqI/HTDKlOTMaJZd3jdjA8eM7NOCLnxoMulKMJLx4O8/fICRZxu1FYu+MNKyu7q8noyWwuipMNLS7xWKDZt0LPqlyB7LEqxXzRavEYM2sHk9QW1ATmCzCzYoNW0VGOQ5FfZilg5b15k6tRz/tX3PyT5ZMjT77GeTR1TTahbyWjPPAR9xn45LDCYbqmXgQ5+r1ejnfg9rvzWqgc8mNUZXnxDzIO0Z4YaRBCONwSYjnfrOPQfX9j3anQLJz2mwNaVbis+QE4b/1f5yLMa7jHJ0oc3Kk1H2YdCt1OZ+vk2kDrKc/fFcCPSQEUKOGMNHMJ0ZkaWa1RXWIy0VbjLMMdnkqcS6yKiWVddlA8CNHOm7jEQburxgjjclI3vdzx89YJRBzcKIVt+kMCsjRV2065yg5T8zsjKHOGcl5LZbTAwzI35vFWmSp14JBCcMXKGwgN7tMyfoA80CyyBYiuNAAyOqtZbAG1XSWhVsPYHLtKtp8os8YtUvGZBDWdXFfDHrwWK+IawuQOCnaNFkRllBygSyXYaA4FRgUaEgLBlLlXKjnfg9jhmlRZb3SjVnAk1GoTwmRk+oRTkpFDWlimB0lUdfGfKItomRv8ZxnRmNDzCiC7Zj5JNdiyx8jBGtOk5K0kkWxmj1fldGFhvY5CkydJwksmcEuhQD1/b9LqNa6JX+f98xKm29y4jjz/c0lECmksnIz4bVGoN5i1FNRb/FSAHYuaBXed4xqnGzbDtP+7q2Ryz62RkMMKja4pQsT6FAYQUaHvRkA6mR6JPFvoGSAoMi008hPLPfRQ2fx8MJRE8YnuFgWpVR5XicHAY28DQpAPE8U/MhZSx+PBhXrDb1qabbwtT0uIv5gu4ze5si3ed/6AfSVxU9mRXmz7t4m5GUe9r1OdD7TVAzoxYsRNdgFGOsMOHTZu9XRloZoTCygqFbRvIBRuOQEdth19oz4qZEIB7eg8qoBaNgxetPjLBj1LGBZ3a0YKSqGG8y6thwfp8Rre0bRhyrwghkdMnvRT+qHHnWRKUwekBHOYqxKIljRnKfkVZGlmF8m5FOjBCMtsLIi+xE0DTObaSBZ7vmKOibnJEai/vieQeuKOUwEy+RjXQaH8LjV7/KN58c3LptRFNb1hU5/W2rLvUglkNNs5ftZ9ELV2ua5W5mukDWbEQXmuCubJD7TI5cMTLKxwcoNnn5QUYeBCuMahruKl9DgaQiTkYa7sU9Rk/BeCC3f3NVCdN4YgTUWBEOGbVkpMko/eiklIxsglqcI1Om9xlpMEIo+WTEq18mRjoxYsUiFe/MyJS8MbJ6g0NGWhltpXcDtwoO7p7BGZ3uMKqulroiHa5UkxGv/TFGkoyQsS7FhkvMNfbJGemeUVoXUAHrrjZ5hoDn0nS0Jkt+SBeIrogDOhwGNV9kQcogmdZf4sZVK0KZ7oFrq2dwdbaI8ub4R9wvLIlJc9vV2bZL+xoanYKZg5B+ey1PjzkHls10bHiJfqPcT7Ujl4UWg1EZYWKkt4w0fUKm4mZGMjFiP4zRAp518McYiSnlG0ZyhxHKe+n5qq/Ct4z8GrEyvc0oysFx2TFqB4x0YqTBaIkJtuE5MhLGqB8w8jJ06rHCqKk9Z8MYNbzHKBeNXMzIyMbsBXP9DtG8x+gUCkmchcUxxjuMaBW1bOvEyCyDmdFIRtgz0uDGMoOmD1BVXOQ7uLisQzsQtQNexh1+kppZ6ZOx6Sd/rfqDXKkxIYzSU9eEW3tGPpfRJ6XY90TF/UUgt7Pzc4AdAW+Cw005r+03nMafwselOVZ9RUYHYvcdr4EFXRhoBBpOYOAJ0+Qxk5I5Z/Wr2btHjCSyJDm4ZDQH0mJ1AN5lxH//CKMhG17b73gYv+643GO03WFkq9LbjPAuIxP6i8tR1qq8xyiPL3Dl1c4HjHLlJaNaC2QyVhltaGpl2Jf2FafhRz1Ge3+E0QYunA0ZrEb8n4zcMrzDyCwRMpprVbit4IaRVkYuR7Jhk5c/wEgQT5LfM5JvAB7QlrYI3IfiYmoKRIr2OWHowIYzdRzsmQWM2FJbIW6dJpGayaeGPfPTI/w4mn2maWX6k6v9CC3LZ5Ruwgq9shrECljDN0sMhmDBhosNvK7QWOEXxMEy7vMqTUG2JXxPMgLg2tkY9YmRFEZ6yEhjRXmL0fgDjFgFea2M9ICR3mP0iuFuxBGjMTFaCqNRGGUcxzg9YGBDR55ALeApYThkRHM+XAeFTY6JESsu6XefLC7E1fINRqrAVc4hQ3bvcctIbxldcU7WQJHNdsBo3THCxEgmRld0vBRGa2EU9mlRhZSjDVewcG8vR2SkdxjhDUaKy3jWdejQ1IZ24cbqyNCANOXN3F70AXVTjJnUGyD0s/jNDVc8IjMoiHtkXMA0Y0TnJ5NPy+fn17mh6VW+4jR+dV+1nPLkK5GteWxjx8CrXc8DW1wNItJdzM7cRCc37TFGYePGfdyj9pVhZqSHjK7Y8Fj82/cYXcHKznpv+3xd8Z2RdFzwDav+Yoz0gJHOjDpe7Co+YY4YyQ0joJrrdxmx7BnXHSP7/j1GV3kKq1KnPldue0bperzNaMMFX3HSX+wamqnaULAw9y8ZnbM/oUi82NCrRI8ZZbYirZF7jDY/g2PPqE+MNBg9oukpP3rISP4Ao4bX1+ex5s45AU++UgBRQFKCMwSyyQsW/RxDyffYZ/q7Xc5g6tINHfC0IZ1geSTY985HIBCeEkIJ6JWu2M0arvKIB/0HW/0CSH5qgP4a06PlqDn3AzkhrZ3WioYlFADfn+IfEXSk9UBGHZu8YtFPH2SUJxOZOJLRCAYzo36HURFs4vEV6SpPeNA/gYcox4HJoFFMRldXHimI9xjRMrhlREElI6YpbdIIHmB7gV7dteWdxgEjM6ubHjHSW0aQ6BFdSGtVpjMrI66mgOIqzzjprzeMOLIzoyUULLyfua17z6imXiujAVoHqTSSER/2tOBTyH5lRPsiGeWZHbeMqpt0zEgOGVkvWlvRmBaMIAoQNzTThbnrvJEV3by6iWX21NASdFF1c2gJc4sm13ATFW565f09u+DmGKO89bo05epTumgCv+J30CWoKU8GUze85GCUwB+1aQJ0sXa3Ix8QVIqOdoz0hhFTafcZqWoJZiKYkBHcPMzSYjJaf4gRnJGq4hVfEZvdiktFjhu4qagVRuMuIxwwiuxEKBDrP4U2Kwpt/LjFgEE26wvHd5RAHWIBTEY6MVJtGNqRblFyep/RiqEDF3y7YcT2zYzcDZzY3GM0uwAzI5OnMTGq1aGKDa9I9wCRYeTnNrwcMOo7Rg3VhT5ilLuTKyP7vQmkidg5XhadRTQo980joNC3oXna8RorKzs2sOEij8iinNnEQSDpRciog7maVtOYzSjVZigTqaT+LvI9NKSUQdlwRtNTKicwNSY7SFIGwS2Z8HnJiIPmoCdGKIxWZ3QpjBjjueIq34Edo7Se2PLxA4yYjj5mxBWC6bSZkdVnWJaAkfOaPqyM8CYjE7RjRtNZDMFI3SSujEaY1ZWRTozIJhnJxKgHIxwy8ld2jBQjMgBSXAKTo5mRvskosx9vMYot4aZVkVv3k5HVxcyMmF26wtLkI85l4X+4w6jtGJXK3ZinMyOoQGRBU9WIWZgSZfdGfJ0CnmKYK3PHFfEsRlX3m9boeH1oisTfLSaT3Z3BMwNEX1aLVoxIHIMypSPQ5oMIXOSbwzVBYUozzbMGeMAsQNAPpLuj9RacyIPjGYT0htF2wGgURqasLvQtfQIlo7S28lyBjzEKLu8wUgUumBnR6voQoxKNv2XUo717RiR0xMhiABssBWqW0vuMuGgxXblnxIwCi4/2jPAGo+GM6Lo2L3a7w4gKFLQI5kzMIaMynZMRSxL6xEhg9zFGIxhZHCcZ5eJHy/gjjNw9KovlDSdzamQFRLKKkMeCZWzBPk2/nFpn+Cc+ee78igXAq3xH0yW1GACmy8xng2tX8Wes5H1qWqrWTTR4BgQMvsCj4wqUw1yH5MagV/nqMYyrB59WzG5HD0HJf6df7RIPDT+dg6shDB9n9GCmtr9jk2ApQiLAxIimqnj/9oyWwsj9yZ27MDPKFN0IhdjxKt88hnHxlWV5l1HEHspKlHUaldSeUQ0SZxn1xEj+Rka6Z4TCCBOjSFtOjMySIKOBjlf5jgf91RktMcbhXt1hZO0LLLNOIiPNp51/jNEnZySA7xK9ZXQFlcsxI3eJhMHNPaN0i6gpbFv9gGrXVbUrcPIPlKdqQUsjNC4gU5BE0bBi4Ipn+TNW/VJ0KaGm2UMzT3yF1fJ6wsyBA6zMmEE08UnC4A1TalH8Ag4W8Cq/YdWf0bAiAzeb96GaXQwEWdk7Yw45KS8xoFwJsWPE4BdN/VtGJ3S8YpPfsejnwiij+EeMoNwoVGsbuLpVRqZoZ0Y0o9dkFP1dobjiVX7DSX/xQO5bjCTale7kfUYyMeLCkYosBbow0gd0nLHJ838SRixvz6zP24ya75F6xW844VfvEQPjW/SCk78qGwa5mZ0BxN1RD3KDgXEcMqJMHjHa8ITuwfPq4qdsvsXIeYa7tmfENtv7lGnRhqWdZM0cKxsl0QkBNxxRY7Xpc0wUmjn0AHvmxilu7m2KAbLGc0uuF275QSq5OltayCL/fugpD0Lls0F3z5SwzzGdKFC5QlVxxRNO+ksMaVV8qRQBmstUQlxZMorNk7BrAEsOGOGAEc8ROINlvTMjrkI5IZORD5sfyCPBaCQD7/sxo/YGI3WX5BEP+stucu4Z1VgBMwtMda+HjHgtu9tejlLhUNQHrl5MxEcArm8yarFBcCmM6oY1Y2RGs1W2/jgjm2RXPOKkv0BjFa4L6MzIpGm7YdSCUZ3gldHqyoYxLhwyylO3yKgVRrRU7jHyw5z2jPxu9xlZW5q0JnaDjCFYIM+Lb1A3tgywtNvEQnHBY0ToVRVWrmrTLwtJqISaf892I9JntmAnBTKjx3Azq+lqiiWCiG36TgaxGq44g5vTRJcIAEXUF3nwR5iL2rK/imiHKSSbHuaTkhGQJc3MUtxjZPtZMrpscZ49Ixwy8tiRmluQjIA8YIeMTncYjQNGVrhjBV4LLniC3jAaEyOe2i3BKLM+wYgr5yRHldEyMeI3B7rvjDRGQ/u7jBSZYdBgNG4Y2XtLUdJ7Rvsgsv25+mlSLF66ws9diaAtlczMiGXfDFAfMcIhI1+gysly9RDfHoysRLzfZdQOGPmnFMeM9IgRYt4oBnrvusInZ42Yp1bzDvnR5qn5LChyke+m5QQ+gzhgVyz6gH2hFfcFtDB18vUsYCHUfbzAx9fFiz64FIvHjuvP7zGKe8EjHvAranS8Zh0Q11mNgBbXQqn5PeU0Meo7RtaPjlewPPoij2hjz6ibKOgpVlzByXuafqpMDN5jlC4jo0X3GfHBTNY/iCnVB/yCCHaVeEwyam4lkFG7ZYS9W1kZtUNGV3n0h9tQEzfn0HyhaOi4YgGfITMzSkvuLUZSGO3laL7WFqu3TTdbYS1jdMKvN4xy6hVGPjFjDJTMEW0/ZiTBagtGY2YEbhU4YsSsZLfxLQzkh+QoLSaRBoGnTtPHqeYUTZpaUMMCm4FX5qMB8PwAaklzAc7e4DU1G4CGFR25G7L6ZBpNhg9lj4Fl4Imr49h1asNLyRHnBiIrl+54wW9+rSwOo3nccAphyj81ZpPfS6PtiBGLpGyAX+HKNBhxJTlBdRRGp5gANNvHDzPySPvkl+8ZnYMRbhhteMHv4Eo2MxJnRNWRf3CX0a0cMYaVJnLHpTCiJRfbydVqCIYz5UEut4zwAUZSGFV3M6t2FSa3c/2B90SBrteQo8qoFUYcr5lR/nyEkbzJiJbt24zYR8ZiZjkqVuPEiJmuHSOrfdG1iZlEDMzUzSXpV2l8uXuNPhvGIIxgDcFl5zcvDc+oxYJ4FD3gB7/a/Vpcp1aduSYUST+NwSMRC/JCfHtwVsFl5ak/kxR2DOArLLrNlaBxlQQDtanxIzgUK44WRrJjVEXTLIVNzn5N23A0DhnhLiNuOMqYziis58q8PaMILt8wYlZAw6fOVdqCxTWGkYzaASM6a/cYpZn+HqPaJyoBfs8iAC9Y9AQqwgz8/QijbcdId4z8kYLIWM0tIwvmHzMy2VtwOmDEOEINHFZXpsZxOIltU9kmL7HgJqNW7iFO/dXjLWSUCQaFWkwHC6BvMBIP+oZV5e0XQVtaW4dyUmLqHH/PQTPz5Yqn8I9a8c1pGlEY/AhVWLCHZagDua2WG3LadJ9UUOX6mh1iNJ0+qlUAUiHwOz6BUE35E2gRfcI/lN4avI5e4LHPZKBFgNOMzPcpGDYAFzyheeowg0wzI7sXj587YuSuhFLx8WfPyMugJ0byg4wsqFctogf8CQALko8YVZeHjOoW75pJ2zMSZ+SPR9jtjzhmNJAl0daLW0a5Sr/PyOVCc7JB8QFGD8HoE/6EdNPuMzILhi3vpW3VdUyLg3JwgaVHbTzLnp7SfpMvYwS3cuaFrH2ckc6yTtcYKtA+tEkINdOnEhfcb0B5wW8QLN7AFJH8N0D/h0EsnvGI8l5qVX5vDrvkhOX12aLaWZ5M5KcZgYHBEd/OwjL+J96P38Fc/Jzmm81CtoApsEZ4oEsmcR1+/gW/oeEECUbVSkpG7DOtjTz7k4wySKVxlT2jnJj3GG1+epOAdQIon75lRCVpjFbUDNE8OjUrQEbLxAhAMAol79c2RjwHJa96zMisnmNGMo0c6w7mdlYLg4zSfdrwClo11aXiZ24ZGXMySjmqfUlGufy8xYgLrdfB4OvEqNYvayxUjE9QUdmJb8ko7dXZRXubUVom6fq/XM9j7biq6GdUjUdTOzfUwPYVgIUvqeUpcgpqudwIxs5zkFd89omxTRow89IojY9jOJBBmTo52I6T/57BR/p7dfKnhWGffsZf8Al/8gG0n44NzVNYnMT26auvKMeMNBh9i76YkfxRRjy2DljxCTyu7y1GmQvnBB87RrbSM4ZCgbfv9R0jvlMrDxVn/BsedozGHUYDVyy+6iajtmOkbzBKNRE7OHdy1F2OlhtGY8coA651kThmdN2NC92QyihbVt0rizr9xRnlhL/HKONZVVHcMrrg+w0j3DBqN4waBBsuWPCABQ/o2ABnxJAB09zVqkgZzZQ2JcVsqwuW09LaigdRcD+Irz6RUrJy4hd8Q8ODrzRmWXQv223eAAb5WJ9QgSywGowrnqfBali8Iz20esYRGBxKv5halM/vSEVR/TdF7nSt16H7sGLBJzSsuIAnHrfIWVuwz8vY/WrN2z8zksLI3JsjRtbPtTDCASNxRldccUZd4XitPSN9h5EFvfrECHcZ5QY5+ARZ8AkSjDx1HCnsW0bLxKjdYfQ9rC4Eo2thVK2fI0afsOHyIUZ03dJCOGZUJ3CcyxKM0vSfGakz+gw71+Ixyq1nRuNAjkYy0j2j7oweXEndZ6RvMnrFhhdXMgyers5oQ2YiZ8u1MkIwOlvrddU1dvthWNpFubnEsLzie9SPp5+e2ozR6GqQUpClNLZhQYcdQba4hTGnVsW12LV0MLU4A4+bn7XAyszspnW0rtz7QVcw9pLXfsFv+Ix/snuUMyV4DJn9oSLUwkickbr/XRlljMfat02MUIRYdgNqR6K9+uppbe2xiYiMaGpWRloYnYN5ZcSiLgYq6TMPzNuXa7p1oDujf3RGZWU+ZDSw4ATVLRjZ+v1cGKHch+N1j1GJwYCVlRs6LsViEvRS5k1z+piRWZhkVIOx83rPYHS6nbmwzYw6rjjjd3z2WNh7jKwtLNI6ZsS2m8LfM0pK9xhxHlWrcma0TfepQXsyuuI5FE6TJs10hUHLFJOZ9ZZKA2iaUAPW+vm6958d4fsWmMr01uKa1SZ8LWqhr7QgzeWyJd47cg1FwViI7fdnEJEuzgDLW5lC5K5Fmo/VW2uW4gwtO8oKBdT9EntGNpG+xqDRv82t7MeM0g82RZCfSSuMO3qrj5yMerTnmFGLz82MEIw0GDGFWIrAUOMa9v4Ro3bAqN0w2vCKb28wwo5R+tgp5LeMuiuM6l6yinRm1HaMzHm4ZZQB9WSUNoG1c/O/jxgBr3icGOkdRnMZt7lwyQhxj3Rf9oyqbCcj9XYbo0/ouPpCk0s5FdSe0SjsFR5cjT1VA10vukKAqKYtQmlm9RqiWss6MngyB4pSG2dQdA78dHAvyQWPOOGn+BQnxTL51zxnYwQE1kQ0tLgqUJWLR39jgGudPM14Dh9jI1ec8ZtHt+GDcA2NXoNRldFlYnR7stVtu44YsUWppGl6dlyx4suOkabJHwNNRmmu5nUro3bIKC2iNEOTkX2Tq+cn/Bqt7ruYQU70rFO54HGSo2rmznKUiokW5/uMLujYcMLnmIYfY9RiEs+MamCPjDIIe8Qoe2Er9wu+4gG/RLtnRghGZGaOyhNkkiO793z1ejfGOfbl5wyKz4wGrlgnRuOQUcYCLzCLi4oOEIU02xpCyAbmBV/dDNb4Ukbiq5nHlBL9QO4PAPjU8B7nNSA+x+90vYaAULiqRaDeia7XIuQZ1TVotCo4WbOkWMs98/XuKHt8r+GT9Vu/FgHOjE/uegW4QlhEf2akbzKiATozUheoFKasaVBYIdBb2YhkdIn2sa33GElhkQ5KCuLMiC6qndb0ot+Qk3qJ+3SkS8Mo/Qu+ginh2dzfM+KmtGSUiuItRhaP6bqhppeTEVkYo01fd/J1xKi/w4ivbz61css9J9+rfkdOajIS9LC40opmrMtadZ+RTIzGjlFzRvUciuYEbPHt2m8YDVTlbYpm05fgVi1haQtWqx6lTrviBb9Hp2dtztRSinquKOAlYVp5AQ2p6gVWK8TusWHTM1Z8RsZDaj6+4QJ7doH4WYTMByxT/ULz+9np07ke2WdzNUf0h0YxtTM/c9a/un9+GxTjSpDKlBmYmZH9vWckoMNHRloE8ZjRyYxkfcGKT8jCnry2MXoyYfKDWqiOZka0orj7Ml+7x4jfpWAyXnDW38I/57inqWvjXhnxEyOY5p6HHI8c+4wJfISRuSSqptDyM5XREhmGPDiGKmT5ICNahRtQzHMSskVnDUYv+nuxVEmAVozJ6iu+FUb4EKO0njK7MzNiBWgyM0ZXZ0TFVGtByOibWe5Re3JF1JjoQLNNWwOqA2f9zXYwlptX3y31EW8312FkUUhmhTN9xdWB2tgHXAUXU0RcIQAAIABJREFUfQQjvlWAr/oMaDX4EnqNUcwBTcYsNBRBBlPz7EpW0dHViICVNpz1N/DEol6uP7QbI1RG7YYRDhnpDSO4oGUxjt2PAmurpwCquOiTM0rTVP11HryCctdbRozZmHB9hBEnGtvLz4gKXvT3uEeOq61gZ/0dc4Cweb/2csTA7tuM9F1Gln246nO0JSamKi76HfkoTgQjREs+wiirnClzyWgF05uRoVDFi369YURL6EW/fpARpX5BWrfispuB22TEyMT1htHQvmO0BKNX/eZ7TDIk0IKRyf7KuXn2YiK1dwN4NcEYS2ioJlyNy+ZKm5qZHbIUFeI1RCcEJ3S11Zb67loi+jxOPyrKohUZNMv4AgUvi3moj6uVQAsg20E/31K3T/gLftJ/gYg9YdpSyFZMxJO0mF3I/s+MbLCOGLGIzMzfPaN0dyhG1qaho4iDRipabhjlfgcmwWZGc9zgbUbjkJHigmf9K77gX+xEAV/dWUzEE8Uo2kmIjKS8PturGlH7WjBIi+yWEZDjOZR87V6XiOi3A0Ycg7TS5rgOf/aMmALfM8q6DAv0XvCsv+En/LMdCQCmR7/tGKX1kleiC8sJmzy5KLK9AGN4ZIRDRkznD6XLztjbE3josx1EnAkNKqmlLdKgw7XcQxkub7humINlVVSpjTlxGqpgdb2EXjYIubEm/cI60bws2RUFc+dc9Xqp4GNk2Pz01P55v/S/La9f253aumsGTamNOZkFDU/4N8DPVaT/XX80GC3QGNi81yiMyFArB73eZcRVPd0zgJF7xCQ4BceZkewY6R1GXKGOGOnEaAlGF2dkE+Y5GOkBI7smhY5ysnfr6sloaR5b1GSoP04TWU25Z1RXXB4/R0YLuKekxXv3GJkzMWfOjhmNwhBvMlJYASAUzuj7ASMtfalWTwZBa8A3rSx/T7fgUhmNA0bm6lzD8rjgyd03ZoeuwYhBVMXAtV90/f385/5f6M+gSU2tnm5Cdgo+/TK2wMgtg1JZN2GFKVtMotT2XJloxjOtZx17xm/FP68BodvIfRb+2AAvvkrzx0zq7kondydmcUrzE7t6CATvKd7TJ/wZihFZCWtDnxjZ0X3V/1+ip3a/dAmSkRfXHDDKSXPLaBRG5EHBuWU0Jka2qmYBXTIavvqSEWsKrmCBUZ8Y0TKwcSSjE76EuMyMMLVvz4hyVF0dHhoDAKq2T/mIUZrxldGGZzxFBkCRmwD+GKM05WdG2c5jRrQwto/JEeZYRVqCe0bbjpF67Q9dULMaPsLIMkl6wEiCEcdkPV8e+8AXv0hNxZgLkH4yg4AbaN6zwam9GPVmXCH9H0WWKFdNmv5/aviODSKs22D+e4CFXXR1KDh0HdJU48Cm6V2DtjQ5mY6ioqIpx0CTmdWPACxv3YQBrrcZWXXpfUZ0x+y9ucCmrhoINWInbKl22F4PsxJuGXFHYi9rkAQj/mTAMvtARpbqy3jF3hqqcSr9T8RI32RUd0u+z2iRU/S7MqK5nhN6vMGIifpkxDak9ZfWUJj0YDxQo05lxWeILDeMrJ8Zt5sZsRBsK+2vjFiflAH0XMQzMDozevW51tFKRuCYkWBdVllPy6f2PP6KL/KPLlipiYiLP4wJZKaEqx98EmSMg+Z3+oCzwqBpRJdkwys6OlbPklz1BQ/4KaAzAJRFLrWOnVPGYyDSMJRnd/KBs3OtP0WCn0G0kK4UU2BAk9X9838MRZiM9IaRTY6OdsAohYwBrQzgpoWQn63BRz5SkIyGvuIBXwoj7kugyU9Gc36I1a+0HGZGGt9HtGcpV+Ak5YYnewBzMvqnEDpG+Tm5KiNxxf/jjCiH9xi9TIxUNbJtefdeJkWuoPkjwYgTlgsIGS3IAsJjRvT7Nz/XpEFkwXNk22ZG1bXLVf2WUd7viNG8Waz2xmTDFO3Vy9wzS6JuzWeBWzLyhMAY2igcZ/0d6T9VeyCNvmpKZxYAMfG5X8QMmsxapAbMtI813iLOL/o1jhjjQ4jsAJ0XZPSbRrgNWC8+XF7T4xuaPmkv/imVGDMZColr0q3hKveqj4gAkRrws371a1RGNTjHcuxUpqyrSOWYVYAZUGPtCa+Rf5PRmYxQGeUKUa+blHL1CrfNx8niMzMjCmMPRjReZ0bsx6s+gg8jskaLZwBqbEGnPu19dLbhlpEcMMrS+MpqZoSJ0VD2tTLq0x/aZtVV6hH7oJLYYhLfMtob8hz7a2Sr6NIrgBf9Fgr6iJGWK+4ZVf6VUcYz7jGyXpz1d/A0d2716HqNeUHllXy4bwVoqkNppDyNv9gDf0OzpslJCyDSdqFNUxs2nDAfZoIYpBxsdtajs3qZtCRdDHtvw0UtUss8dvWp2A4OYh00g7iiFo2xnekq5eAzuNX1ipfxFfNx91kr8DT+GsfrJSOAIaXKjCtXK4ogt6/XQi9F7n6sJ20no1gJtTI6YdMrrmqPiRzoE6MMyFFoRtxvDqIykJzK4C1Gg4xKP9PaBJ71N2e0xApNwa7BTv4cM6pxH/j9uYv2ltGmr2DZv5RHCxqjF1z1BTTXZzmq7iuVHBVAppGTUd2VyXbQ0qxydMHL+LZjlDG+txhZW/aMWjCSG0Yc30z13zDSFZu+gPGUphlwXnDCRc8xF8mI92Uf1tYWGcrU2gln/R0/4Z+QfmT1o4dPi/R282zEkodHRrRrjGBM8AVXfcZAxyLlcBIxqwLi1Wd6xUWfscon0IPkasAt5fyp1671F3Q/MmKSVXFVkQyoa30/9Ug/xWrEEuCGBS/6O77gn9F2jFjqU3/ES26PGWU70mydGV30GXrACDtGV33GcsBIg5EURrmC56SYn+2aikV2jAZe1PeJqILbxcmIE/AFXz/EyNRTZeTxmFB2mUTkDy1Nmv4XfbTxEt8irwMqMjHqegUUWOThA4wy5lUZoTDijo29VQm/7qs+FkYsq67uhhWu/YR/vplrWRyH0p5bRrUtGaNCKI3K6FU9riSeTNABiJi1KoIFJ2x6gSqwyCnGMWNKHcv/8D//9//rL/9y+gIgDqq96jm0nfn/87kC6VtTkDJwmP6S+bGxizUG2xVFffbobrWp1YR5hHpH7tGfC0Z4jczUzP5gBmsYcZiVBK/zqt8taGgyZvcVtfSo+IG6/kCmq54j+5KMMoI+M0pFlkJjyqEykgNGuMNIdowyq8HjDuvKecvI3n+fEcrYxSSQlofL7hgpNM723FyO3mIE7OVICiO3zKTBHhc4764UCC44777/HqOsVmVoMdsyZ6/m+FQyErzH6DtElsJozIw0Je+qL3cYobQLeItR8+8mI+sx28wKXwAHjNqOEfcXZWBVpOH8m762BSfTwMpIt13grL+bL6MEtZQLz0U21SfOhqjX4mddO827V32Kh7vSXBqaufaufFhu2YGqwIvyGZTzTsL4DIA0B+up4ogBoJOSK6ZpYYvZWHUirzcwALVzFe24dC2McMCo3TBi/IaZIbpuZLGVPR1pkanHAwY0GC0ei7GfcchoeFCWPvh9Rsmquky3jDQYXaMiUeL5FLeMtMiRTowylXfMSONeyciWn02vZcrkomR91TuMFMOtCW4TN0Ydr/pUGKXrlYwyRnPEiAvintHmjBoWfz5HkVVnxKP9WmF91q/oqIxqooGxuMpIdowGNq0V0FkoZnt5sm9kRBtk6OaMqLjT/Y85oorWmrSuG2zHxTL5UHRJTHPR9GEOulb5cTWvOfST6zcWemh8loNJWEOH+5jlWQouUNaxLQJ7XNErRISWtUFPtyQ3w9T4SQ282io48Dq+F22eT9piGfEWCqEVRuYzWtAzC7t0xygHX24Y5futtG0J35GrMJ992rCWgT1iZKb0pi/IQDRiQqbaZHUf08/3GQFwRk+HjGRixKpZY7TAnt1iApsbv44ZtdIeY7QcMOI9N7VHGvBw2VtG2T9j1AsjW8gy/lAZUTp5olW7wwgTo6EdF2dE2c9q4mTUlSXjwxl9AlTwMr6HHNE+T0aY5KhmdhZkapgLBJWUxSj4rBeDQkbxEOdg1IKRWRiVkUBEsDZZ0bwghaCH37DhhPP4ii/yT5jNxWpS0/fPNFItcq658w0vMOPtFN2OKlBVN2PnCD43nIXAqCWjVnyO11Jh1c1v1XTMNBLKatE9Ws1V2dd6ZMpqQSvfH9p3jAz88/gdP8k/xTRLRVo3BtFc5QqVocdkNJzRAvrVrGnBISO7wp7R0A7FJWr57VrpUdPNSd9YPsCo3WUkN4xqWtz6YXL0j+8yqulISMz6YGThw3NMelPpZKTOaD467pbR4sr/ApSNVTXxWDNjQHVb03Ulow0XXPW5MGKcpcFS6PVE+D2jDaxfOo/fg9GcSOBYLRARMMaYjHLUxJMBV5ibrMGoBWe6YpmKpUpLRraXpMiZNjSErrfLWOlqzU40nMdfA04tiqFQpcZnOkhLE2ySXPU56vaHr4RDO8AnIgEYenWNp9NnI1rsDw1ShWvNsvpNwo5oDwWh/lhmoUemJV0poK40NcOiE6NrYWSC8Dx+2zGSNxjVI9qS0UWfItMy1Gr4jRHcH90zMv/aGHlQSuFxkOGrb9ah7BXCMSN6vP5oAOVZC4rcZ+AWQTkte2bErfWWwqTpbq7e24xqnIByccvIJ5D2+APXKwqa1u8zGtqx6eUuI32DEQOzVhP0fMBIAnPG8m7lyBjlAU60VPfJheCmZGT9P2b0GLE1ytBwN5plCcmIblplJM7oIVPPQ7SJNNGAXX1PM9HNzBOcx+/+aLWGrtyMssYRYply5ZO1BHx8+2WcQ8A2fS0dqwGkNPWYkuQ1eT818rEyXfQlBs4Ui/oDUTICroD7c942FbzqM57Gb7BH5Y10f9TcJIucS0xKPlKPM2HBQ2HUffu84jy+ev/JSHeMmHV6QPifCog2vI5n0LTfdP+g4Qw27Rl1P+KPcQF1AaW1ddUX6CEj40Ffd9MNFkNaPT70hOfxeypz/1tUnJEdPU/hS0YSjDhmqt12M+vAeXw7ZlTc0mCke0Z0hfQOI8apuLmqMjIFpjeMRsgk62nICJWRIuSC1uXL+L5jhB2ja1y3MhKfF5XRUH+ur3a8jO+gm/omI3kw96IwehmPLudkhA8wWt0ahbu0bqx4SGBoR5erNE4ias263ZirLFf2x/GvseJT+9hq5ykoVzB2AK5p1quercH+pLDmE43BnK6bPz8C4JPVGTCskxX+t8VhTEjNT3QtGoOv0+rPg1Gg4sFExWVwl10GuKi00j+VGCApjGwNJCOdGAGC7/1foRMjOejTzOiiPLODjE43jHg+aLW8eD0EI6SV7L8P3XAZT8Gx+t08WCcfyygeTFRcx3NkexgoTUZLMGPQLN3LLGKqJn0yAh77n53RkoxKf4MRktGru4t85updRoqZUUxUFPmxKURGm17xOp6tnweM6lGByWhMGTFmt2rMZmZUHydxxEiCkWLgsf/bm4yGB5Mp22RkiswUgyn++p0ejGh5MXCfjBCLcjISvL689CZ+keECzC9YNWWPC9LqeB6/haayBucJPCOizuIR1XMBl8EwVisyWDigGT3mw1AoOCH9rAbNjI0VgT3gOs6+eqgLR8YW7Fqm/FQHnoc9M6TpGoIHn2+3gjXCZSL0hA0PHHWkUjNGT+O36LO6qVgZ0bztuuE6zhHseouRQsNCiThN+PP8cVcqHt7TsPhJ0Vc926rBaUC/2YOlZDS04zy++sQkoxI0LKuo/bs7o+GMuil/zoEbRubicBw4XvcYmbJ7Bt1iMsKOUZZvJ0e6xXtGoUx9Iq/4hIYFV331lZVKy+MkrriS0Ybz+HbIKBe1PaMeE3y4pXWfkY3d8/jd+uULYzCiQvRe2aL5XPrfgi1jOwzQ8zMMplNxTYyi4jQt2U+fviyt+kWMRxjQrD83IaS2WvC9/zkunBWLNtnVTfurvoQZx0lvAZMq4PRQGUHO7AF9wlBMcA3o16JCse+vuPhBOVzvu5tgrWjYl/EtosdZtJUFSYCZzxlXIFgyqFV4NRtUGTVn9K9lzZgZcYJYVWFmcNIC2TOyg074WzJSZ1SyQqFA0oQUmFKklUdTnPEpMhra8frDjJDKDFlaHMryhhFitXzs/wp7UPR9Rhev1dgzmuJMihDq+H5RDLMcddCfj0C9W5+izRiJK3mXWZkYbXgd3ydGIxhljcTMiBOzylH/EKPv/c8QydQnYJmJam1c9PkuI3G55PL6IUaxqJQ9Kn2zvSHWjAcwIGTarfmAmYZsuoQfZwP95+gotTFdgIueozH1WlaQAruGUiCsY+FzK5B7H4q5pWXVVa6qLcxxQXNzfnFF8+DBnYGuG57HX0G3hA+95f2Y1koNjhgIWwlM2y9+YAlXAfF+jQNGgOCp/1sIARmx5s8Yubk7MVoPGGU/2L5RLKBk1N5g5HGeURmtseJ1veI8fj9kxPhNZURNSKuTn1uUjLawvjQYSWFkfX/sfwlGY2JksaVQ1r4CJyO3Rt1c5lix7iXjBPAxyjGbGWHHCLgMPpdkZrTpBefx1Rl15AOmGajHHUY9GIk2tBtG1YU3RhqMBp76XydGQ0dYA6+Rrk1LBqrBqLqnozDqO0aTXGP1fo14LrFIQ8OQmLCMBOfOTmqeuaaCD+l56n8pppStVK/jO0SlaKryE/4gN8XUQqXceQlk5SPNbSo105xuFsYqb3lxC6Y+h4+5eDT3RfkAoDTjMy7tJa9+PUbXrV1r+fxw85iB3Cw8kgNGqz+A5rH/mwsEB8xNWDUr7ZhRpn5vrRMEI/77mJFObQp/2QPOsS1dHmw/jPIBQLeMLEg5M+oTI2ZPRqyyGXykFN0yOuEzBK3IkRRGX321rA/rdnlUxk98c5feMsLEyC2x4t4kIxRGCxoeANWw+hQajF71MRhxra7XOGaEHSNuYmRMkJZ8/pkZ2fkXT+OvO0Yd5/E7FnkAC9KOGPFIB7qslOlklD/JiNXEEv0CFC32hqjFKcQ1P7UztS9rEagFGYj7PlkYtk+kau7MKlRNz1WT0XdqebEHCquUNmh0nv6exQ3U2wJfkRD3fh32hKhtXMw3DsDDldrVv299Yy38ggc08QN03I8MwbzDiK/dMhpRAFMZbXqJ7cDcaTszcsvE/4g2LHcZaWE0c8snZCUjOCOzMJ4AbdjGq8UotAFhIZAR4p7GyCZTE6aykxEmRqvHc/aMbGEYzmhQRrDgcVRGr8bIr9EmRloYtVCui7uabC/HNhZCtyBmOWplZc8+08q+jDOgMjFK6zs/j8KokVFJ9+sBI4uZZTzjbUbW/8eRluo2XrHiS4z5PUYhB2AxVvcYi3i7dbKo5YiRKX5pNetBzUQtC1h5CfP+rEjbcHF/V7HKJ3zv/4rreAnz1jTXvP8itakpCFaGMa3J+21gRSmDVBmsI2wFS4SpEbnvfo22n8c3PI/fbODBXbPifWIJtnlzBNzdhIS3lTGKPNdxzyj3XiQjpojJCFjlAd/7n3Edtg8gV7f5mmntYGJ0jTThzEgmRtmmI0ZA7rgkS2P0uzNiPKYyQmGEMGFN5ycjvWHEzMAxI76+6Wu4kQ2VER8fICFTyQiF0TIxqiw2jyWkHDHm40E9Zgim9dgZiacpVW4Y7WMze0Z06fi6h9YLo7otgfOM2ZcB3DBiNa6g6RqMuGmO8s6RmBmRn+4Y2f36ASM9YKQ6IAI0UfP6OGE2zw+nedsjECb+xYbVTyBicE7cl6ul2hI+KM12ouPj+Jiy40YqRudjpQDTQxKCucpDCDSvzc7yCVWqitfxPSLITCVxmtctzDXyzsfO0/y1mjX6fbJjlIf79ImRaeVF1rBYeN3z+LZj5EFE7YeMeCLzzKg5I+63SbPxlpEGIwaSN3+AjJVwfwtfPwXLflowYnZiuBidQgbIaBwyugQjxgR6UaZDbSdtE7uOXbc7o3qS2Z5Ri4m6uRxRRiwwx3SisUpGnOTmGqzyyWSHGYjKKLZqd7zsGWndrOjBZfU4m7vxyYjWWGWEuOfm2Rd4z8ISc0Zdu7sZzkge7GTw8T37ybkQRWyVUTmrZGKUCYJagRvu2o6RuSJAa7IIA3INK1Z5QJMHL1DKg3VzYiEmlGUYHtG04SRf8Nj/4iu0bY4SN1cZnLNBNHNr+l140raVM7M2oU0aziBQeCMjMQ12w+bnCJzki/9uRUc0OaMc2N2GRR7AoBD9ukxz2WeaZCQ7GZ2CUTtgNJzR0OFFNgtW+YSn/lc38y8+ZCxAq4xMoW16deWAOEKPbhMltvkKOIpSfp/RK17GI07ys60w4XIwoIqolBWszsiF3DlURs0Z2XutMFrdlM56gRo7MDkyhchCpBUPeOq/BaOclJWRu7DKOhpP1fokgQKLfHIrEWHGV0YWLBwQccunjD8ZvY4nPIidT9vhwUhkwDDcGCx2hIC/zqtkSlkwxxXIyI4hjGKtsH5Y1ZyMqCQWnNBwwnO3YrCZUZlr3j65w0jVvIKQC093s8grHv/gCgUCtDHmBwWbnwLXuoQ4wrei92PR4deEoAMnfLaVwf0kgoQLVB9Z8GWd5qG1acKF2qa/5iuedSazH1mMxCiv/n+cvWeQZcd15/nPvPe+V7a7qr0D0GiHhic8SBiKFAmSA4qkSEorrYaalUazkpYTG6uRtCNObCh23IeN/bIbsTsj7UxI2p2RNHKkSBmSEimQEkkYwrtGw7ZBu+py79Wz997M3A/HZN6qaoCaRjCaaHRV3fe7mSfP+R+TqPwYI0epP7HYgXPQ0QMhb0leiPMlxK2M1lpeGMW7xCh7V0a+wUjuaRjrYkeg8WVSx0BfG8MLswkjdVP51KZ6kbCBkVVG4GsV4gaI2Qqg8iOMPV0pKN2HlKeX+z/jhk4ZxUUWQxUD0TmIUeyBEEYcaoX4LJLRSUOmyo+QJYJ4jhYzytlbuRKjwIyiF4IgoSN7nUFCYTbMuima6yjN6JR+iLHv8yYl78V5GvWYpmijiCzrSAyPazKC6CaOvR0p1JMsX1xHCAHOb2RU+7EyIqpFrBhOGBlhFOK9JzLhPDLiQFueMyBhFNeR91LMxf6htbLZI6w6cVXiYg2cXSDLOBKjANnftJhsyND3SxyPclm4oY0TU15WqynlYaPBgm5Kwyc1uYReNYEYm1odaOVCRZkQ02LbzWGSKWBMRmXPibstBiaA0l30WUncJJeSvS0TpyFtYBRC41mgjOjnDNmjWM8IwaLnllCHEp5TxpYNbpoWlNg3qtdAnK8Zs0EuyNRwp7zkuQwsYGjp1qHE2A8R74vNIyOIhpBUIiaM3AZGsTdSBU+IK+351KshhU2REdYx6nLj10ZG/QYj9y6MiJN4OhLOxloKHqvImyiGgvxchlZGHcYoPU2UElEQsOrNic7S0IfYm5Cq4Q2MAjYwkpSz22wdgbzHJqMi+Zyy6Q16bpHTxWJgcmYkY/PidQ5ivCSMBB94KSP53YP2LTHgA1+zDghskXhAKMfFOmSDT08Dg7EfQOdqhvTkoJ5+iwwDt6LGwAcHY2LbtzEWNMqejIFDTXXs/KLlBcTGMZ98VHLlXKjYhSPXWEaYee5xqMOY1WuvlZYVv+g0TpS40wcH50ttD5fT23meTbgZI6TiLzs6vFnHvo+ctYr1jGSA7dCvqoDsUkYmgzGZMg7sWjpuIpPwRhwMaRwToyIZJmEkHsnId2FhNOyQMEee2YUaVSjXMTKbMKIGKCijCo4ZCVcNqfgYUEaIIdLY95Cjre+o4YFwWnTou8yIv6cyyjdnxEN6LW+2yIjXEd2IBOmBiYz4YmO/poyCMuLsBL/7mhnFzyuGlxjVfryRURBGUWdLQ0VaA7KpxWO0GPk15GhDsoBimCIjMCN5hxWHzTRYyRq5f4cY1YFupCeDspGRDw4yQUuqR12okJnC5DbjMfohwBoLIFd30xou1krq4l0oYQL0xG0XW7Fv/jjK4Zs4u3aRPhgccpNh4DqYzni0WiC32qNWF16sfaaVZ1DD4BKxSqydGhJI2WtAK5+Bz2rsnjgIA49R2cXK8CKCl3yyZRNDU4AqP0ZhKb/fzmcw2ZrBdGsrMhMwKFexMlhA7VmhNwWCkUH0MZ6V+YjEyFJMD4Miz1G6ErWngitjogoPGBibY7KYwUx7Hu28QFX3sDq8iOBy3bRxLD0gntV6Rtq0l+WAq9TTiIxid3Arn8XeuSNY7j2NhX6LwxtqRabFYGBNC5PFFky2tmCymIAJHv3xKrqjVT3NNAwwLIaJa2py8AtVVzazbVjUKD0Jk9bkrN4HIDjSCazBXGs/Zlrb0M4KjKoOOsNFDOohmzu5SzZg5LqYnzyCQztvxbb2FF6/+F1cGqzAcBO+9JFksMjzaezachgtv4JTq2eiB2g4Be7peYp8BnvmDmE8OIWL/WVIhW9u2pFRqNnIQNdhBmrddqj0vcsvOchoBKIwMpyOZ0L0zaAJA1DYkpkCOTMKzKj0ffX6bLKOJFtCE8xJ2xi5NUxn29TbiZOumows/9y4/2SvxZDf+0q7ckXYhgnIg5O4K6jbBP6QIQCeFWdjLEaO3KHMtrF9y1HctPcBHN1+E7ZObMHlhW/g/3vh9/WbhxBQZDPYte16TPseTq9eSGI8IF51SBAdAxMgpMQGfRmSvQACptq7cXDHzTi4/XrsmN6N2fYWWCMZEoe3L/4l/vDlL/FpbfVnABaT7W24bve9OLL9VuyY3ovZ9mzja0+d/3N86ZU/56/g2NtYMjDGo3Klfj4VD43BzQd/HHftvhZ/9NSvY6UEwHMHimwK++ZvxJGd78H+rddifnIHWlkB0bCH4wv4o+//OlbLiThnEwYwFnnWQvAlai+lx44zLAYz04fwsRt+EucvfBnfffsFiJcDkDe2e+txHNt9O67dfhyz7Wmcv7ADv//yH6sxMSbD9pkjOLrrDlwzfx22T+/GVDGlb8T7ER595d/jsQsv6sIRETO3E7AGKN04xr6GvcZsGg8e/yfYm13C7z3/nxCUkUcC/za5AAAgAElEQVS7mMfB7bfimu03YM/sAcxNbEdu4/tZXHkCf/Dsb2LkY78CYLF72z14+PrPYfvEDAws9kxk+JOXvwJtJzcZ5qauxrE9d+LIjpuwbWoe/bUT+L2n/j3At78bWBibY+fMdbhh7z3KZWHhEfz+i39I4qFp66b3XFAlcx2skYIv8mSdrxEMUNgJuFAjSxiJgY+rO+g6otF5yeh+XkeSlTMgcXnoOpqN8HwokfYh+5Gb20Q7Q0DPLfLhHC+CkubINHSlvZbzv7PQqXpdUO8tlq8HjEZjlxtjTEjcn3iHotg9+lX6IbZMXYPr99yP63ffjT3TO+H9AOc6ZzDVmsXqmDsJTYGdW4/iht3vxbFdt2GuPYPlpb/Bmyt/oh8ycEwkterGZMhNpkDZYmlNPJ3gbezbfjNu3Pc+XLvtMHJjMBxfwpmVZ/FU5010xl3k+Tbcf+Sz2DGzT09psuQ5Duy4Hbcd+CAOzR9BbgwGowt4e+VZPNM9g854FXm+Aw8c/TR2TO+hEx1eP88NBz6Oe695P7a2JvHcG7+Db5z6Li8eACbHnUd+BvdddSd8dQHGE7eZiatx0/4HcfOeezHXnkHwY5zvnMQzC9/F0mARtXc4tPch3LTjMLa22nh7uIiZbDsMLOZmr8N7Dz+Ma+cPohy9if/y/X+HgaMF44PHtq234KM3/hTm2xO4KG8qAFunD+Lo7jtwZNet2DE1D1ev4e3uGUy1jmN1vADnaxTFVhzf8yBu3Xc/DszuBeCx0juF1y58CxfWzmDsamyZvg4PHvoQtk3OQ4RYHxyKfBvuOfwZ3LLnNrStw188/a/waucyYQgGWTGPD9/0eRzfdgDLy4ss3lns2Hodbtn/ARzfdTMmshxltYqzKyfw0ttfRWe0Bm8M7jr0U9g1tR9tm6PvSvK0kOG6A5/ER45+HKPBq3j87ALuvuoBLPbOwcKi3d6Oa3e+B8d23YH9W/YCocKlzimM2nMYjBdRs2CwZfoADu+8HUd23Yrd0zvg/RAXuucx1TqMldEF9OpF5GYCov6nBwx5axLmUU+HRQ5jyOU3njIvwkj2TayApHUkYrhHvCQrGiE5zKhWaOi6GjoYzlDIdYPi4UgoLAatDjS6v1cvYzqbI2/E8BQ17UMJZCQMlwSYwE4h65NG9BVOyQYWb1GhX3eRhxCCxEdiMMTTkGGyZRgizwr8/Hv/LSxqLHRew7de+RJeWXgOW7c9iJ+YP4IzK2dwdO8P475rP4Vtk9Pwro/V0RpCaxqvLz6HtXoJM9kOZCbDwd0P4O6r78YTr/wHnFpbhXSukmGQZ4mVZZlp4bajn8O9+2+Bcz2cWfgenj33DZztvI3KczeeyXDt/k9hS6uFp089ChcC5qb24+CO9+DWqz6AXZPzqOsuTl36Np4/922c6pxG5Su07Qx8qHHdNT+B6dziifPfA5Bhy+Q+HNp5B27cdz92T21FZ7iEYKaRW+kmBfJ8Cx44/o9x2+7rYYzB2cXHsFrnOHrVj+EfHPkQWhZY7L6Ovz31Hbyy8Cw65RqJucai3T6A9x7bh97aMzi9NkIrn8P2uaO4dd9Hcd3Oo/B1D5WrkFvp2aEXvnfn+/CR45/BbFHAuw5euXQC7fY+PHTjz2L/7DwMaix03sC3T38RL156HLt3PYyr5w/hXOcibjjwcdx36FOYb7UwGC/g2dNfwksXnsDCYBGlH3NtyBR+aM9HkYU+nr3wOOrgsG/rDbh25224Zd/9mMo9euUQkxOzyAzUIE9OXY2Hb/lFHJjehhAcTlx8DLBTuO+6X8Sde44BYYyzy4/jpQuP4s2l19GvexCvcde2B7BzagtOv/11LJcjTLZ34uCO23Hj3gdxcG4fLi09iq++9gg+ftsvYzh4E+eGHh+99Zdwzdx+ZAZY7Z3Fk2/8MU5eeha+fRQ/dccxXFg9hQM77sUd13wYe2a2wcBhqfsWHn31r3Fy4XnMb38An5i7Gm+vnsZN+z+JW/fejb9++TfRGS3TRjSxuQ5GUvgV14XkkAlXLjj4MELLTiuLzBT8PThLIZtTfxn9PehmpUzSMHB61EjqnJsqAwnVAOsoRm5uo5CYQpgCdRij71YxbbdpRq0OpYaKoiVJqGI07A3wQebZxJoRFyqMfR+TxZTJJY0DQF0W+hhklWSuoAkGz57+Cl6++D0s9BdQB7pb9I5dd8LA4J5j/z2m21vQH17Ck69/BS9cegIH9v0YHrp6Eq8vnUJuJoDWDH7oup/B8R1H0O+fwqCqGkZCXDaKi+nfxTW/3HkDz1Wn8cKFR3Gxf04jLFX+s2144NoPAa4Hlx/AZ27/CPZvvRotC/THXTx/+o/w1NuPYnW0RrURJgNQYeR6mGxfi/uueT983YWdOIJP3f4p7J3dj8J49MoOnn7z9+Cm7sAdrRwvXnwGBhaz04fxoes/h4NbdmB1vIq5VhsnFk7i7mM/h/cduBvd3kl89fUv4q2VU6i958Ii8KTqgOuv+jh2tifxxsoq7j/+T3Bw23HMTcxiWK5icfUFPHvhVfzQ8c/i1KUnMHQemZ3CdQc+ggcOPYiqXEGdbcely08in70Fnzz2KcwXBifP/TWeP/84FvqXMHQ9ABZHdt0BEyzee/wXMd2aQX94Ed85+TU8f/FJ9Kohe1GO0msBmN92G27acQhr/ZO4Zu+n8eCOG7BrejeCH6M/uoBHXvs6Dl/1GbTqE3h9dREBGfZuvwcPXf/jmLUVBq5GUV/AmV6Jj9zyP+HY/AGcW/wevvn6H2Kxv4oAKVwDhS52Cvcd+iRaKNGtW3j41l/BNXNHMJUX6JcdvHr+z/GNk3+Oa6/5aexsT8H5q/CRG/8RxmUX5xafwHNnv4fzaxdUZ7ph/03IDXDkwMO4qT2H8XgFr537Bl648BSW+suoWCS+befNMMHinmO/iOn2LDq9t+B9UlcQJBSSDIrTjIg3MofVAMag9iOUvq/XVaQDaXhxq5nwCOz8+8Ze83AY+zX9HoG9omDEy6cSba1EDhIQcX0SLIWumIBDjZ5bwmy2E8HEPSRhR9BMUYgHtJErQGOfmONrODSlTe6MdNiJtSNFdOz7nPIxqH2Nb77+ZXXHjLEw+S4cmb8agEVVXsZfvfo7ePny86h8gDE57t9+Ezq917A4LnHDVZ/Ag4c+hmnr8fLpP8UTZx7F2MnsSaejzNXyBjKkohCfvvgI3gw1Bn4VhZlAhozLVen5W+1d2Fq0Ye0E7jz4USx2X8czb/0x3lw6gYXeeYx9qS6fxKQZWnCmhmlvxWyeITNzuOOaD+Fy9w08/daf4PTyqzi/dhq2fQ1+7r0/gfOL38DFUY1j+x/G+w9/BBNmgK+/+L9j376fxtZt07jv+s9jtjWN1879Gb726lcwdKnHBA6rKAbdMXsAgMG1ux/EYHwZp5eewN9dfhanV19Drxrih278F2ijh+fPPY3Z6UO498gncGTb1Th/+Xt4+tJFPHzTZzA3dxs+ueuDGI3O4mvP/S7eXD0PFyoMfIcY5ftxZH4vYIDx6Bz+9sRf4OTSCYzcWEU3TbNxLDs7tR+FMchnjuGOiX04v/IKvnXmK3hr+QTWxgPs3flhvH92Dk++8ruw+Xbcc+0ncef+u1COTuMrL3wZP3zr/4B2No9P3vYraJkxnnj1t/Dts98CtCkv6MJFCLDZNOYm5xGQ45arP4bO4CxOnvsrnLz8JC6tXSCRFMBy7y30yluw1HkZL134Ht5YPgH4KTouDKf/TRuHtx+hk9EP8djJv8CJS89j5GRyNm1il23Hwfl9gDEoxxfxnZP/Ea8svozKS5zvOURYxyh4LsKzAGJ4kps2XKhQ870eklWwhtOOMNyYZhobVw9JQ8WNOaf9WfbUEFAckbQSVYyYhEwODmDBUnSMnlvGdDafMJKrDln/o0WpoZMInvS8Y8pWmTaFMz7A/K+/9fOrM1eFrV4h0C8axxYrJ+tQIWN46lbZWbz/2GfRWX0aL1x6Hi7E2YGt1hF8/v3/EqPemxjbOeyemsfCytP45sn/glPdc5jNd0JEVfogUgIce/KtiYVDdSgxcMv8ArkwjLMGIurtmbsebTPG5bUzGFSlUo6DWunvSbpVfBMHj11zx7Aly7G4dg7DutS6ECDgmn2fwKev/xjeuPhdTMxch/0zO7Gw8jS++vL/iwuDFRw78Am8d/+d6A/P4aVz38DJpbcgAaBY/Vj7SENaJ9q7cdWW/egOzmNlsJKk1QCb78J/975/hWl3GW+tdXF05w2wfg1PvfElPHnuabQnrsIHjn8a01nAuaXn8dzbj2FQV6hDib5bVqE4y+bxwes+i0uL38OJyyfgeIFIuX16QZMwyrIZXDN/HK5exYXuKdSeU7uckvzwrf8at+/cgxMXvo8DO+/C1qLAa+e/gb95/Svo1xnee93ncO2WnVjqvopnzz6Cs71zEAHOIuMydi6T5jTm/OxhbGtPYHHtNDpjToFD7hTl951oXfGZHWaznZDBRpmdwnuufRjZ+DRevPA8xp4vBjJSMUybYBg8Pnz8v8Xy8hN4ceElVCFeJB2NQsVt2bkamThFXv6ebGrJFFY0Bdu0SY8zIo4W/OzN+0NpjcsoPNEf7CaMVPZGFB5/MEYBHjPZTk2XZhpSJRdX6bshRmUYssBaqCbSO2tXzb/67V/sTO/3W0i9p41e+SF5DrBcxurVSEjxR0wHRYuXIecfCLQmrsMv3PfP0UaFy9038MyZv8SLCyfgAim+pR9gS7EHsZeiEJNIm8YQOB/ozs6B67DlbYZK8QWKSRWByTYA81Kg1K+R3LZ8ZXS92nY6Lm5eEHt3fQCfuemzyOGw3DuFZ898Dc9cfBJOOh5NIbYZYPEpXIFRenmL1JzE0W3stWXz+OydX8ChLTsxHK/g9OUn8eTpb6EzHidPHCNfHxzdWeG6mra7EqNovPwVGMmiz3QjREY17jz2efzwwXvh3QAXVk7gyVNfxenOeW4NsMw2cAg7iIarsY5iwdZ6RnKiNhnFcuh0IjlAPShb8l309byO0vqedB1RK0BPb+X6r2NE68YluoHkPWL9T4bCTCg7OVyl/ynoevAJI0PP9Y6M5MihtZxmoWRgz3pGgb2k2XwnJHWbm5ZKDusZVVzmnjIyMBiea3fMv/6dz3em9tVbBAhVHcYLb7Rs1Vi1fjRoI6jVE40hdhDS35uZ2AmLCoOyi9JX+t/EKtahwpZ8N6QzhUIRLn5iD4A8ihUUdgLSUyBuM0LUOESJFlc/xIAxSWdJkTDUwko6CSFAuvuoDoNb8bknY3ZiOywchuUa1uqVaPnZ9kpoJrn2IAU7nMGwV2BkjNEFEg1KjlYxi8m8hUG1jCJsRVSspRoxZTTGwK2isBP6OeUzSxzaZCQusBQIxb9PizFlJOXJVDdgbI6Z9lbkARiUfTj+bHGCGK2koe9yeXIU89Yz8nyib8YopspjwlIZhYDM5pzap8NrS777HRlVYYQhh2dXZiSFUu/GSE5uifWbjMSDyG1LD0NJP4sxBQyGrsO1GiH5vH9fRjFJGxnRfydx3KtXsSXfhbCBUTRmZRhyX1WTUYBH/2yrk33wR+/+QjZTt4FAhoIflFJIbO0g7zs2uMgvmWCs7hnijWRl3UfpqvgCILc+04fLTI6h76BtZ9hmyvg2elFVGGPgVmKxClIhllViPv2tsZxadJxHlq7JEE9sNlKxGzG2ZYuhIGs/1BZgazIgeIzrPsb1CH3XYaVcrLJBZpJLbE1oMArvwCjwE0i4I4Kth4f3JUZ1H95ThR4xkoUqpfgULg7c6jsz4s9qTaaMxDuUDR6v6IuMxCUXRtTZ6DCqeujVHS5B9kloR5to5LvrGNkNjFjB24QR/Uksk6d/aB0G3cjRONEaGPm1KzKKbvVGRqnXKevJigctaVJmJGMB6Gvp52fs+qedvwB7e2GsHrMYCfnvQ9/h+Re8p1TfaDJKDQDpd2kRWBxxIIy0lN2YBiNjDEa+jwk7g/QqClEsSj/A0HevuI7qXl5aazJDpcdd/uJMX0AAdKMTgFqrx0QIEnfVsSWPE5Rk+GoNaeyxyUkjm6IwbXTrBf0zUZNdqNGrlxoPL5kPESjlmcjFMPz0LbW+shA1RRSoMk+9iWRzSBu1RYEMuTYSSa2AgcXQdfUZaGHl6xgFSKl0nAngGox0GAtC5BhqWuJXYJSZFrr1ghoTqV51oUKvXuaiGuhmsusYaRlxkDdcJBmnwAsvdnbmMj8yNPUBaVCiRZ7rVLKU0cB1NjACfzaRN2kjVQ1G0tkrg4wiI9EDNltHUeHPTIFufVkPJWFUhxL9euWKjEKII/CbjGSGZhRGdSJ8CMhlkrlkPhCziT44zWpQg17kY2AwcKtqhFJGqcGhdVRBBNKYwYvj79R7ShjJAZTJ/R/KiD4zMYoNg+R1UbpVBNYmI+5l8SHYEBwGrosCE1QxxkafasOb3XV6Z4JYwxBgeSKRdlZCWrxZW+BWYhIrqW8j8MaWKTw5WuhUF+NLhldDEecfeMR+f46j+eemTVSy8eNEI494dZ1Y7vj9JE0VZypw1VoAj4enfwaug8JM0jNJWivENvqUkZZmS9gkE7mQJ0Y4TmuOjLLNGQXa4J3qUjQWXICTS8lxEO5iuIWRYdHYJIx4viMzkq+JhWwSE8dUotS/yF0X8melH+oCHbhVtOzUBkYmYWSEkSkajEyyjsTz8vrerK49Y8hg6Vh/ZUTvsFNdhjTQ+VCroUgZhU0ZFQkjFgm5c5pqKby+s8gjg7Tqb2REXokPDpUfq4c2cB207DRyTsOGDYwQP69exs1Gm6eZ6awVIFnbBtDrG806RmhMhu8mjOpQYVCvMiPi6D1NzZIGRQAw1iB734/c/GvFbGjLSRN0w/FDI7rLgd0iUYqj+BOzKGqxQJ2lloWSRuebiVOqxJhnpkC/XkVmcvTdKgrNWcvEav7OpjnrInox0f3LkOtiSyvkZOR8fE7b+FxiRGCiIFeHkj4Hi5FeGcXvExkF/V61qumZPmMMRDYTyhJGJsbp0emkE0gYDbgcWBjFXMt6RtjASFKBwsua+P5E6FWXfx0js46ReAnEiBvOrsBIPAxZZzULqU1GaZmx4Q0RGfkGo2aVsWS7Bq7zjozwAzMSoy+MRIAXRnG9x3fP3qqGX7l6CVUY64kvGZxwBUbye8pI/GRhbBuM6oSRk42mbJJPDmOMeslD7oehAzZlhAajqpuNbX/Qq63JqWVctYWMN3lQD0IEw4xHjgkYgheH4gTtYotTlQA+MZLQBkGMDF/DBhJaFsZvNowIPTQNU5GadbHmskSoRp6sqMRt8j3TJiDLcySldl+6QGM7cGyQE69j5Hs04HYDIwvp6ExnIggjizgDUhaflwWVPDsJX+sY6feMjOLwV4OF8Vv6QoWRlclcDUbpfZ9eGaWLqsko+69iNPRdGofHVYcpoyxhJHMR4jqyDW5xXgeiQPxujPhgEkbygS6P30oOOzmQNmdkGozAjPJNGGW6N/Qgg+HnjcZT3oeKm6Bej9rToVNzYZiIo5IFSRmFTRiJQfL8nCpYKyO3jpHMh5EDPHocPjgslqeRHvRyaG9gBAdrrLF5kVtpWpFxeRnHUNIijsSAyLAVcv/ITcs5dShj5ERdlQUo48TJXbPJYvXqutV+jH69gswU6NXLGkJEg0ReQaoPkGtJm0osdB0qfSlixaMWkpbxej2xRDhK5wyIICTDVYauu45RbHqLqVjRCmLRDbmHwkbcXR6gEsBDfdczSgftyMQui8pTbJmZHP16WU9wNQjBr2MUV0Fawlv7khnlrF8Io9ivkCmjulGnIG68ZIqGXLgDGAzdGk3IQk4NhzqDwbAnmuopkp5MGeW8eQoxE7RxA3dLBmmmirNE6Xl44C0MC77UW9FTRlHsbTJK5rEoI3riyo/fgZGLZd/BKbPNGXFTmKWLvEd+DQWvI1lLV2IUEka01q0aKmEkxsrqOiIPREYZiCcYm9touM/Q0ayVPo+SiIxCwsjpOwAAKwtzUHdgQCKJ8zW8T2+aipZfT9XEBZLYV+5WFIsrszzFIoqVk6o3VeJZNyGtgDZUp7qkC10WbWBjQ/F/Ae/5ghc+/QJkchLVLMhUpniCZHC+ip/AtODWp3T5BBvUXTTCrGAwrEkEFkY00SjemSILbyMj02Bk3okRosfQZFSz65ixEc/RKS/y6RWFVTHIuCIjGj4jtQX0WTYy0tZ+UygjGc4SGa3qohZBceTWeA2kjJyGH01G2SaM5LJiA5niVqcDcNkoyLamSek848TXGLo1iDdmYNEtLyEOd3KNdYRA68VtwijnEfvvxCj1xpqM5OAJxMgUyshvyqiKmkjCKD2A1Pvhv1fLlDNlVDOjOJ9CvleOFmQEgvM1Rr7HjGhdd6qFBiPxDkn/oCxL7apgY3wI9F2HXoYxgJGpPlG1l1MsikMBtafhtXJCyuaKlpseWQZxyMKpGW7lS/TqZcjU6yAeDTJ0q8s6VCW6RiKWOtUEyJ2XOYuO+y8kDRZvWkrvN1VLm6SK6WsKDN0aRBCj04OqST0Chm6NXoYRj4IZhTislwyKTxiV2sBDjExklMTClsMXWTiR0Qi9egXUetxk1Kkuq3BJA3C5NkKEQKxnlOgUzChbxyhAagbYQ1FG0cUeuC6QfI38fBcchq63jhHXvYQ4cYwYyfQqzwNjmowoxPRJ5sYkIQCdljV3Y5Z+hD5nGaJ/QN+jW1/WTAqto7zBKBp222BkfgBGflNGxHro19R4pIxqX2Hk+8pIqpJDAOTKAAnzfcKo8mPdV6nHcSVGJO5T12gAMPbDhBH07yMA3XpRGcn8VNofGZx3sDaXXlSgMBNAAEa+B5nSLLlyxylTWag5TxkWL0BSTOI9qDoLcp2kDTaKZOT+1aHC0HUh9xTYIGIXNFxYqxYharGB1ZOBXlQUg2I6iIyGWOMUiAiz8tLIXWymh0dujV3PmNEQU98yEwgh0C1QmzCKqSsKzYhRDM/ktJEYVDID+j9AF4kYcGK0ljCKZdqWha/NGUnYkTISV9dqiCnuufyS0Czd/OLdCcchzznN+ORJNZgCEwjBNRhlWnMhjHyDEYVnLd0UxIiFP2YjIS8QZ0JKKFf5sTICG24dBccDcdeqRTb+1DAlU8fES6Lf/TpGVhlBTTo07KCNJYySA4i9UDrRs4YuY2BQmAk4TxWuwjYycsngJ2gHK31dO66R9HvKvNt1jOTgDgGo/Rgj14POxg1A1mAE9OolZRSUEXkrxgRYgyzQA8c5FkO3pt8oXZRpKsgk/6QqueR+RUVtTtmStFWNOlToV3Qtm2w4EZS8r3WQaW5aWKsXUYcxJNWYxmOpiBNdOLKbLjhUbpS4jFY/U+0rDT1ErBz7vj4/kOgMiEq8nDZD1+PN0mREl92kjOymjEKDUTRIos04zjAIo0wZUUiSMiKdZ1EFWJswiqc61OAoo5AyqiGXUoMN2npGmcnJhaYjkBnl+gxanMQCpJZWNxjJZTd+AyMxAJK6lMMllsKDD6PIqPJjDocsF+LFsM3D8+145BmsKSPhHrhKFesYyToicd/5GqUbMXOZ9UCblRjFW9IlC6Nfryc9h4X87jM2NmMu946McvYccvUmhJH8Ul0EUddLGZEhcfx+S1R+hEHdSRgRa7kNPhpRi169xCMu49q0yBA8QvbAj7znC2ZmPCEv0/CCrDhuRPKgUtkn5c3pPyLIGXZdRAQSV1v+nlhKqjrkQhn2FHQQK6h3Pz0Rx05GjBn9WTK9yHHJr0TC4j2QSiyuO708mueYxr30p2M3gGF3M4SAYLj334iVje4leLRcHcZqCEWhd9q7Eiv2IqNoNAy3qmvJsbG6OeS6vAGLqsLIb2AU43jAcE2/CKgmYQTQ9quVEUy8b0OU/8jINzinjCTUEQ9IZofG1C9vDq72lVBKGPlA1aK0tkRglJ8dh8eIZhIgPTqev2dkVIdSRdXNGJEbzZ+JPbmR77NmE70FSR1T0UDKSKac2yswsusYOYxcn934yEhS+H4TRj441TsCDIfQ8R2kjJCsQzYtyV6w+pnlMMhMjiqUGLseVySTIdnIKAqbtI4GelDSqzPwvaK0YmWlwAQhnqhSfSZ1FxZR8ZXUkFpCE60rQtLIA+jitshQe9oEksM2sJrn1So9RFGVNnChNQZiQOKdB/S8uSn4lAiNZ5TnTjtqxQCKjlL5ET9nnJsoVYlpIY78uwkyI8Dw15q4CDYwsldghGQR8KI0wojcatnowsgkjBzodm4NhfjqvH5Nw4QANO6FyDj9HHsOan02YhRH8cdT3iij0vFaSAulgIRRHMsv31vmblZsVKWDuMkoS9hkqkvFzRwSRrFvovIjjFxPD4zIKKn2lBJ+FulSRhIy5Cw+ygYmRmn/xTsxChsYqWe0jpEUva1nlJtWQ9SVKerUBeoajIzJ+F3LZ27W+EhzgzAq/Qhj12eNxujPE0ZhA6MCMvNTGJFnTZk/S15MjO2duLj8ssl9iYtWBSSBEeIJQotAsgt8JX2Sr6/8GL16iQyJl7SgFADR95Z4XPsRRHjksEPiqnjjVYDUD+hGZ7Gq9pVadvl8YgQE9qBeA/hnSwow3iQWL8aJsb0wkv6JAsO6+66M6ASh2Ru1MuLJ2yFWnZKYuUwb84qMEsMF9qKCVLMarNXLAMCiIZdNazVfzGgBpsEIEH1HGBKvQS29HlmDkaT4hE9qjEnhd/p3RAtSQ41sU0byNXKtZXpzPTHyKFnwBQxCwsizbpMycusYyXg5WYeVL3V9mCQEUaMOg9qXyTryGxghgBkVykj0Bvn88j1TRjX/bKmwHblek1GIFwJFRnWDEZsASFUqZTWov2lQr/LekwuhpOw+g1RcR0bcRKe39wVeh1TWEOBh8yw36hojQ27b7KbRi8lMCwO3RvGZjN/nTawNWhL3IcCC+gZqvnFL8sEkQvX4w0AzI+mpLBtCbkSPJ5icji0UZhLL1XwSAjUAACAASURBVAUVV0lJLyFpLxEVyb2SFy6KPNRdrUOFXrWihiEg9rfQBpKTRbyu9YwKZWRNzlmSoFWrwkgCoPRuDEnvyp0XIu7RaTmApLGEUdjAKGO9JDIS8S03LRSmjZXyAqSI3QfHE6J8wog2t00mMakinzBaS0rKhREZtVLDk5QRlNGEnqIivlKWRBhxefV6Ruy6y9fKgUDPQFmPsR/E72vkekKZyRGrDq0ygjIiHayNzLSxUl6ENE46ZuR1HcXGNpm3omtJRUReR+v6c0Q4F0YU9+cJI0q5FnYSegEQP+PI9dcxQpMRJHyAfq0UjuUsgI79EGO+NErYp+FkkxFfdgVhRP+vMLTGV6uLLPJmsC65SUpELdpQUAOAAC3iSIulojWjLS7xJA3KoUItUn2HGNQdtagcnSkIEyycj+q0hBpi42mTk+ssH2SlPK/eTBziAcit2rGKkA2bFpjQ76XjqkxfygdlYY83DxscqdWQlvZoTCIjMIshnwxalAP6PGl6LmZynGowzlco3QADruMQHUQWeBBGIWUkQrIwEg2hVoO7UtKcCcnu6OMqoxB/TsJI0nOiUVSeBwnxh1ZBkq3f5oxK5gL9TD54XkeREd6VkUxqqzB2AwxrnmOaMKKK4NBg5IIMyo0vKWVk+Z+V8iIcqEVAMmDKKDQZeUQvUDxfYtRSIRKkDTcYifFZ334gWoVsVllv5GEUmzMyWdyHGxiVGLk+RnVvIyPvVcCVbJnTvRYxpWlty5nF1fISGbwso65Tz+IcpQErngthOdYjd6Vfr0CUaNEBxH3xSVwJQEMZD0ehjPQAhPSSnJCIUqJNSHeedFeyRfSxo4+s8gT69Qrkqj6Jg3PbYhlTNpFHjIut1lGoZU08HBrVHu/qkO8rJ0o6Vo3ET2JEFYv0wkgzCJCilsjINRjRZ6r19BSNQk5MqbdAyogr/q7MSL4f341hJ7gatskoswUzCmpMm4wyrqOg7bueEQzekZEYndhSbdk9p5OyX3f00EkzCZsyYuNXh1I1CiveqTKKlzenjLRSdgPzjBlRlWmvWtFNI7USxCgRpvmdCA8LYkTDZyIjNRKAfhYgekpyYAm/5oVXGYu1HgPRVVRTtLANRljHKKPBNa6v7xIpI8RQUw7YdB2ljFyyjkTQ7o6WvfXBB4nF6KXI5TMsUqrnQXdnjHwfIkbKLdni6oqABQDGWCq4qpaRxkf0Myp9QLF8VKwy5ot0PVrFPLZPzeuHiCXVcdCMgUW3WlBBK7cTaOftuAHsBOan6JIjsZYj30O7tRX7th7GlvYM5P7IwB6D807dzqiAUypKXDVhJKGJxJAGFrltYeT73HRWJxWDdOpOT27D7tkDaNmcGY3Rq1cSPoZfFFcZJoxy00Irb/MCCPo87WIrds1eg+1T2xuMAi//br2Mdk6j7qW+RE7N2tfqSUhc3q87EFFUdJLIqIT3bFx4SpPcXi7CKnkRtIAlQ6YFVyZHbgq+f1Y6OuPdnnEdRXGwdCP0+cBJ/7xOxiWIUcpMTqd8iIVN4mTHdZToBxyOdasF3Yjai6Lp0Rrx/g3anP16BRLqEAUuFoPnG8vYEBrDxqlWT0C8tMgoqHGVvWBNrh29wkhOe+9r/bvyWcbsmYqYLqGlXiSNGGo2GCFlZDdlZGAQHEKuSmugyUgyjdDzaUMjuDwv9Ktw456b8fr5b2CttIBp4Y5j/xBXZ+fxxZe/jumJ3Ti6507sLPr46smv08bM57Bv2424ed89ePGN38bZfuA7Kmt9cHIL6WEdDK6/5jP46LGHsRXL+D+//euYm78de1o1Hjv7PTh4zEwfwefu+SV89dFfxemhhW1vwT1XP4wb9t2O+WIN//c3/w127noAH7nhE9jWbuE/f/t/RjVxBDftfx8ObjsI40cY1jX2bdmO//R3/wLnB0NMTu7FjXtvw8XLj+FcbxUeBrcf/hxunB7jPz/3B7ztpPCJe0KDhzE5rt55N/ZPT+Dps3+L0gGT7b340Tv/R7x68j/gpc4qDu26HTfvvxe7Z+YxHHdh8y3IRi/jNx7/LYz8ANfsuA8Ht8zhmTPfxNAFTLT34lN3/jO89ur/hScvn8Ls5AEc23M3bjtwPw7Nz+H/+No/xbh1ALdd9UFcv/tmtFCjXw6we+4o/uzRX8DzKzRTYsv0Ady4736858D92D0xwr/75r9F33NLteo5gSsZSRsYuz51/MqkKFlMgdKQmWlpiOe95+YsuqQGiR9BKcig2otoDggyLMdg5PqYzLckYQdnroyInx4jP0DpB2hZKogT99+abMM60toKPhWl0cqHgNy2aOkHGRsY619IQyvQrRYx19oDqTKOxikkGz5g5HoorFzIFL+HehHMSG5ulyxLzOxYWCOV0MLIKCMq0qIq5ZEbYCrfwp+TMn2SfYmM+ij9iAsrJTciKef1jOJdr1q+bgw8gFwqooOUDST3BxmY7L6Hb/21fNZPxKlBGv2rpSQAOT507GO47dp/gOWlx3FuNMZDt/xTPHjwDrx05hFcd+Qn8MOH3oe52YPA+C08dfF5HN73EH76vb+CA1PbcXTPjXjs1S/CF7vxwRv/Meb8ZVwcdOLP4aq4Gw7+N7hvzy6cXhtiwvSxd89DuHP/nTi6dRseP/M4du+4F//wnl/GvD+Hl7oD/NR7/xfcuus4Lq0+gzeWl7B/ehb57K148KqjeHnhFLa3A6bn78Zd+47i9KXH8cjJP8QTb/0NLo0zHJ3bjvO9Pu468mk8fMPHcWDbzRiuvYi3+0O8/8afxw8fuR+vnP1r7N37EKbdBSwMu9FQMKN9uz+AH7n+4zi241q8ePa7aE0dxk/e+6s40C7x/Ysn8GN3/zNsKzxeOPNX+NbJr+CZM9/Flvnb4Yan4dt78YlbPo+7DtyGozuO4oUz30Q2eQg/ce+v4ch0gafOv4hP3P3reN+BO1CNL+CJM0/h2I5r4SYO4uPX/wguLz2LR078Hv7uzb/EK8sXccf+W/Da4mncduhH8enbfgE37TyOTu9VvLRwBlfPzGJU7MG+VsBCv8MniHSVBmS2QK9apvGF8JCWJgp/ZMPE9UCbBBq20eJMRrUBjXVEU9DoQNI5HgDGbkCLHOu6aJGRUOf6WmwltRYirAPS0xNPQNEFpE4iQw5q1eZMAIdZscaEvla0hEG9hslsFjIhrcHIFFirltCyk0izSpERP4MaTpNwkWs3k1mrPwCjgIBSGaU7lPyZsRvwheA/KCO5i0eGb8v8FS6vF34JI2MyuG4xzN7/ibu+YGfKdhO21MrLBzEwxmBhbHDj9p14ZXkFH7vl59BffRazWw5h++xB9FefwZ8+97vYvv1OXFz8Pm498jm8Z+du/NVzv4GnF5dwfGsbF912fOrmn8TS5b/F9y88h9LFOxbBS2VteBbPnHscx/Y/hNyv4IUzf4lBtg9LS49h284P4gNXvwdvLJ/C/q2HcGDLbjzy4m/ir1/9U7y+9BqOXvUwDs/tw6XLT+CvXv4ytm+/CzNZhZff/hoeOflVvLVyGiM3RgBwZN/7cdWWXSgs8PrF7+D7507g8PYDeOHiq/jwLT+PbPQmsok92LnlWrj+STx57nm4NOxgRsPRRbjWVcjHb6JqX4ePXfcQ3rj0AvbNHcL+uYP47on/B3/3xnewPOzAB8CjwF1HHsJUlsHVy3jsjT/FQj2JqfptdPOD+OSNP4o3Lz2DffOHsX/uMJ567bfxFy//AV659BJ27rof79l9HEvLT+PLz/1HvLxwAv16iNrX2L/zXty4/SDaeQtvX34Sf/f6l/HoG1/Fa0uv4fBVD+PY/FVYWH4Sj5/7HhBaiOIgDWzt1x1MZDPxJOHTW/4enWix2Ivc7jTYicNr001rOVUpGpGsJ9qgpPPQ/bNtqlLlRVqFEYb1GjJLHoPhsEc0MeiKCXrix1qawOFj7L2RrJUXA8AbhdZ2LFCDAUZugIlsijeT6FPUOyWMwrsyCpAZpOJN0OaPBW9NRtCvSfeEbOrKlyhsK3oVnB4duh7s34eRiVcTSojdGCi8CSMLC/TbpfnCb/5sJ9vV30I/RK5Xs/qgUm3ng8Pe3R/EP7rtx7Gw+gq+8+oX8ery29i+5Sq0/BirwwFKX+OzD/5v2IVFPPbGl/Dk20+hDgb79/8IfvbWT+DkuUfwrdf+DJcGXf2e4jKlk41lLoKFhbGT+NF7/yWOThd46e2/wbdf/zqGmMLVW/fhUudNvSjHmhxbpvdiPDoHhGl1o4d1F5ktdCFJWlM8GTkJts3fiZ+5+2exuvYGHnvtS3jp8pvYvuVatHwfF3sL6v6RKyyl8eS+PnjrL+HOnXvw+sVH8bev/SW6tcW+rfux1D2FXjWEDx5tO4nctqiZp15By07qZ7z/5l/Gg/sO482FR/GNV76I5TLgqrlrsNo7g864D0kNzk7uRzv0sDyiWak1q/rkLlL5riy2+FmB6andQLWEfkU3sbtQYTbfrowGdRf5OkakM1T6/6nJqKaLg9lFlbUhNSi+wSidtRCzB6JNyHtWwS4EtOwkcltg7Afo16sNRrKhJYUoGzWuI69/pgOOjNwrankTJ4wMpSCEURz9H/U4YmSYUQe5bSeM5BpBYSTT2moUtk0iITOiqVdR75Bb7+WZ1WDBJxcJrWdEBZMtO4nMFhi7Pk/dmlRdoskI+vWbMgKlaSIjMXzcHwS+8DoAmS1Qnp9YNb/2Gz+zmu8ebI0uiIgg0rUYy2HpG8mV9hlyW6DibsHCttGrVlDYdgKCK9WM4doN+RW7GsUg0eWyRfKwccisuMCUXqMXTPA432xz1Nx6HkBFO3Ot3Sj9iGNgq59LCoECeFQ/rTu15BLPB8p/aepKRKg0/SWMxPPalJHJUYYSgV2/ft1Zx4iLYQzehREVvuWWRq1JVuYHZmRyLeIhRmNi5AbIbKGbupE5QHRXEaCfcSOj2G8i7nQ6y1XiYiBylpMuA3UGV2Gsi3dQdxNGQX8mraNiU0YiRte+RGHbkAFImzFKu2ffiVHlS8y1dmPkejqpW7Is0nhGpzFfY/GujGQYcrw7xACQ+0XS6xc2ZeTHWkY/cn2d3p0yorUu1dHCSC55jiI1MZKRgCmjGGEEZhLgUJ6fXKVybz49pEzUAJr+k7SRdB/KcBxJmYogsjg6qwIK7T/ZUFKY45IMSmz+InGTKzcDkHZPimsXY+KMc910okrlm/M8vIZTZ4WdwOLobUhKiyrpeG5BEA2mRV164HgxBEiRk6S1ZNKXD15dSsnCiHCmWrIwgmkyYtfSB4el8fmEUfycMSYXRi5hJHUBSd+K5vF/EEZkgOuQMDI5CtPmd1ZAFfhktgNABV7a9Zn0HqQDduRuTBHl6FdkpIuZ2dK7knkRsXgtA9VzrIwvMqPmaD9pgBJGPmFEJ7aDpARjtWbMoMkcTXK734kRlFFmClweneGrIaii2aLgOhuvf4ZAov07MZLaGBExY8ZCGPFBLoxCnKkhfyc3BUauj051GdJTJIzos0tTXMwwEaP4PE1GpsFIBE9hJM2TFhmKvGWtNZmRGEc616QISlI48qElBys2C4HmcQ7qDqayrSjdiAHG9A39zjXtyPnyFXIrdWirus1pWSx9dcH1/gjQBSFijICil1Dw6D2L2pdo2QmsVcs6gKX2dGWfhWWjxD0o9ABwvAg1j88nk+SZZeKi/DdJN2XI1QDI5ljPqPYlhiycUfGO1U0KNkuSViRG7YRRrJ6U0y+mR4nDRkZx1kHae5JzDw2lHUu07CS61SJ9dl9r9am42mmVLoIM/ZHLgWWtxDka0g8hhVWMFhkK7bKUDSWeoPydivsYJrIZVJ76JDIe8bcZo9xGRrIBJSNDp6Fp/FNI89i7MmpFRp4YdUpKqzpPncA6NhF0oIonBj4wNjBCZCTCpVHvhN5tzvNa0sbL2id3AQMo/RClG6Ftp5TfuzMyCaM43CmuI6O/ZxsYZcrIe0+z3Ah6zPfmtqUbT+YbSNWYZZcYsKhCRflvW1CcZahcNRVT6M8NAqTL0+t/p5LaWDSSjjKXGLIOdP2b1c0V+M8rOi0g1xHQ55Bcc2YKLkpaIRcsaeoK7JRJbR6ddEVMR/F/if+LirL8t4ZxCsniCKHBqPQlBo4YyaIcub5a/ciIqzU3ZRRP6DgPIo4FpJ8vjGJdRvRSmrlzqlkgI5fbNvoVM0JseGuWkQujlvITDikrKUALCJSJMIVuUrn+MpayCyMqcyehrlCvZuQGmzBK7hIJQVOcOoxJioqUEXcBMyM5/JqMXCyMSmp5+vUqctuiJkXbRq9ebTAyDUaRQZ4csDF0jQOk5Hd5J5nJOeVJGpEctOsZlX6IEYeMUgQ59pGRakgbGPmEUVxhUpsk4SalzyvyniTSSNZR7epgjWW12FPsIi+g9OOGyyuWpvIjmEAnQb+iqTs2xIEzmckxdkM+wQ3NSOABODQLo4wzBpBrQRctNdpwhWlTXprjKc/j68DQvXfIEd0/ee5eRRcSeS8DVAx7GIuQYh/HJeI+OATveR5lRa3UAZDZk5mUHQdx4wKCnEj8AoQRmJHc7aCM3AjDusOMrDKyIEY0n9TQZ1BGdYORTTwX+fcmIy5m4vF19CzRtQ/KiPSVXkWT06UBywSLwraxVi1BhtNIC4DbhBG51fQ8yog9D1mcGxixK5ymyIVR6SjrYZExA/ncVj3VyCgWM9V+zGFxDglJxc2WytnCtJGj0Opf52W6O+d89D3TPrLI4HzNjCY0dDDBIkcLvWpZGUmxonQlr2eUc/GbsBDvLPDPbTIarWPk1jEaYlT3aY/wzBHpDRJPVRmxofG+ppL7BqOiwcgoo5bO6pAiQk1lB+5rscZYa61Rt55zyQYGhW3riUuuU8buUgsuOPSrDj8YAMRpU9LkJCW0cUoyuV8yWch7ujmsDjWp00HuvZBTlUt4gwc0Fkxbfiv1DkKg7lFpv5WyYlL0KaxaHl+k8CoJuaitvYXCtlUUknr8WqoKOS9PKiidEusZWXkJ7GYqo7qjLmLKSDy1fr0KF2QilTDKlJHMfaQFGGckCiPyxljbMLbxkiWbYZRRoKwHhyw6XBkGjo3ryvgipdAajFrspbVZxZf3AmYU9DORom43WUexIEg2dW5aqH3Ns07lNIxl5JK1GtRd1kMK1R0Mx92RkdcBR5FRiOso0X+kPFyqGaUSMmVUsPseS9FjR+zK+JKe3MQ5NhYSoyxhROtI1m46yrDBiEc0REZFwqjCoI5zRUmfYU2Nh+YM6rXIyNPPo3Z2HrrMWp2UcQsj0dmipwg2xusZSXcrV5lRl2g8HSq2Sp7FF7FIlR+jX3e4Dz/mocmSiihqkds2hm4Njjv59A6NILMgeHAKn8jiAjZH0NF4MO/JpRejJe6cGJ+R68WYEFRDaPj0QyLKdqvFGIOF2JTjWPOQ7ytzGGVUOwLFtTLIRRjVyohvR/PEqHQj3pgtSJeh00UQ1H3NuU+F2rFlNHxkJFkP4SEbUhiJofDBw/s4RUxa9IVRZgoMXY/DCJvwixkvmU3ZrZbYtAkj8vgiIzbXyijO5xBGso5ccMpI5oE6fodjN+TBNYVuJlnwogOIzjVQRumApiYjNBg1Rxki2byGD7hUIG4wsi3dmGQshBHH9CZDt1zijRuvMYzrqJUwyhuMQjCa1Wow4s8mhkv6n8ZugJHrIzZKxgNdJsSJxjR0PW34i3NnAel2TuedNhnJjJJ1jCBKBmuONjOWJgnFZpUYf8YxXVI0UgWxcpQqzK3URvClJ2zNMlvoKU8t15JRqSHCYNC/L8NQJV8fO1Izm+vfCZAGGt7urNb2eMI0nRrU+SixvuH0rmUxNTcFOuVl3QQ+0GQknXNoMoUU3bDA35uKfiIjOlXSiUkAFc8MXY+fscko/cy5LWJLsRsgKujCiD6pNHbJSYsNjAr9ng6xyShl1K9WIR2V0qUojGzCSOLtTrWoQhsxcg1GSBjJu5WFaBJG4mlGRhRGVH6MkevrM9Ilx5TylcIgy6KceG9jHb7j9VQURirqJYw0J54wimXt0sMCzox4HlewOaOM13RklKFbXob2T7GGEBmtHyIkXh+glaMNRhLm89xXGJQ8rkDWjHgdIsjKpK3cFMj5QuzKj/X5U0a0h6UplIYVNxkZXgMJo8RLtcbCOxcsjzRRjQABcbYjCj05na+xOr5IsJJZCgJMvsbCagYiNy1kyDCuB9Ar4oIMKMniqcgKsgvU4ESpI9IcPG8gE8g99z7ozx5WPfUEdEaEj1cn0nM4yJwFcYeXxuf1yjsZOuu8Q/BOf65FzmlDmbGxnpFNGAVV+FfLSzEtyGFPykiEwJpHwEvmY+yGzKilP1N0H7L4Tq8eiIyQMKxhlRHFvwgBg2otGmWeNeK4EUlidGGUZg+Wx+f5HVGeH4E6f5uMMgnCmVHxjowQaABSp7zMayOyo3VtGlcRUmNfpYNqSzcCAvh6xHiNXzwdnV5jgWD4d2Ek93vQxCz5O8Soy3E9tamvZ1T7iq/GkCHL9Kwr4wvKSDJAxEgmo1tdB0Bg/6Ngj1Pa6mWv5aqPlfUA3XJRGekaklT/OkbeV9o7IxEBvYemEyB7w/mK109kFGWA5E4UHy/v6o263o5dFSQLkGYb5NZqGIrrevUK9Q1wqEGxk5y6vuHmyKkkQ1ECQjImTuoieAMHqLUTt1FCErKIsZkH7NEAVC8vHYw1p/3kw0pYIBaVm38h7mJh2rg8OoPSjyjuBhX8VByK0eenWZseNBbOqtdh44loYobDhYqrDicgwqi8ZGEk3Z6qT5hMFxQV2vQ0TGimX2PlacpIQiphFNYxGrkBV2bmmhqNd6nEYh5tveZaEsuGcWF4GpUvlRGYEf0Mi8wW78jIrmNU+RKDuquMRFtoMpIuVa+aF3iTuVDT4BsujKKw0MhebNQLXYkRxChyGfiw7pPWgBw0JLm6AqMsYUTryJocl4dnUKVT25iRXM5FjMgzrdmTi96P0cydpOZLzgyljMSYil4RO3nXMTIFal9i7IeQJrBYrEifQ0IPqdPYyIgPSJMy6mGiNWltO2sZEY4y24Ix0jpd6v96lZS65iyc0AYFuBYDOb8gF6sM1QMyKOwkDCzWymVayDIHwliu/feQKtHMxpvJna91A8BYFbT6dRchALktyFqCpzUlsZjEwVWoCCpo7JrlVNhEPou1aoWfMEPGQp6IPVGYMlpSGxllMIbc6crTHZb9BiM6veTil0w8DU5vuQYjo4wAQ8+U3LdBbnqRMLLstpNL67hASMRFqZno113Wa1oxxYwo1kqBl9nAiGea2hYzWoYK16alXchSB7CeUQA1pUlIRzd7VSj9SAVWcqH5ch5mlBZpeXhlJM9IP2MKPgT0qtUGIwtK90t4GRmRIXI8+ay5joiRiL0uiAdq1TBHRhkbhFibI8J4O5/BWrnChjzjcJeeJTKikLSwE5qyzHkdBZC35XyFsR9hWIu2tJ5RiDNUwzpGaqAN2tmUJiBgbMIoQ25bGiaZhBGYkRgs0diIUUdEfhnyZ9RjcL5C7eRmsRq9agUt29bNLy6fTEWqfDytnHfkifhaZ1ZQsw40XhIY4kZXrlQhKyCgdGN96ZLyAcAzJjO6s4INmix+ToRBCkvooGF7yXX5cvzIJCUEGse+PDqv8yIzLoiSUySEONNA0pGREYtSvkK/ohJuhJhx96FW70xK4tczEkGrwQgW47qv8S8xGqubHIInRhBGUpQjoYHFgIVDvQ7PUGo7hmJ8g7dQCtiEEfiEaTISz0yuFEwZAYbT1p5d3XiRFPWftOnNBKk/qNWwl8woIDKqfY1YTk/rQIRomeIlcXzpR3pwheCYkVe9Koq/zKjurmMko+1i3Y2c5gzrHRgZLI8u6M1iUliXMgo+WUeeBGkNB0DjAkf1GnLL65c1MhcqFYFLnamaMqo4y2G44A0ouB2+dMOG1lH6EcsIlPIVRuleI2GZnruv2TMLY6yxPtAgOQEvanPtK3TLJf3/ZDwcKhdvjqp5ATXixxBV7bEbwnun7qJUxvWrFY63uASZYymJYU2QElluK+a4qV+tQuaDOl/zsFXPl/9Ar4LT9BG/+MqVuvGMGkZ6IS07iZXxJYhgV/uS0nBGJiqL62objOTvrlXL/P/lvlRhFHWTBiNjdcCPDDihClNhRJV2/WoVNmQajtReRtdJ7YTVmhAau0fpuF61qt9DGIXgUVi6REoZBaeMDMwVGSEEFHYCq+UlSHhRc2hi1zFK6x2kQrByY/SqFWUj+kHlR2oIxJCqnmUyfgZS7ks/UuNDqUbSLPpVBzZYjb8jI565wZcNiStvkSF4T3UUdkIZiYdU8KFIf1br14k4W7sS0vbQZATktoXVcgESMsstdMoIcc5mxuUEIqiWboR+1WGPmn6mDw4l30AGyCg8vwmj0GBU+xJSP+G9x6DqKiMTDO/ZmHWSi70k+2hZ91urVigUApXFO1/DWgvj0GxqGvuhFjhR2pBcLItMT3SpN5DYLbX+svG0fZebiWSykUGGbrWoKRytl0BAZuMdEJbjqTrUmq6VNKi4/AQyjjPTmB5xxqfoAKT2Wv1d3DprciyOzvH1cHSW1L4kK0+HSiN+jYw6yog+9+aMRK1fnykQ15U2HL2wdIpYt1pSRpLOoo3Pg1T4FCBGpJkUdkKzGikjOV2EUZwpYZSRPCc2YWSQYWl0TocZi8egJ2HCKARKA47dgE+nli5sSQ9L3L85o7TpLKbJSan3WncCAN1qucFIDrWCFzppcRmHlhV63MiXKaMWJB0vG1Mzc0ka0Qeq9yEvhDSCJiN69pRRSBmZVHOgg4rmbQ5ijZBufpksZxqMRONoMkrTvGSIHMsB0qawVq8kelL8rIWd0JBSpprVXJXdshO81wqu6sxga3a/BZLj0KPN/fyZoQYVmUIEkMWH1uHz0NngIY1V8cNEi2hg2bOgTVvYCSrxNXIhTYD0V8QXwkNQ2J2SX+pOGkvlxGqkNOPrtAAADV1JREFUaOMXtq0xajONFxuKvKdY2QWHlm0jNwV5GBLPJS6uFBOJYaPQY5WHoEiItRkj2lQ5e0Mq6IFiY3nhkZHRlHPGC5ny7HL7WpzOnOoPFpZKgVkBJ085YZTUDlBcTYYkFhbFVLGB4WpQ0YyE0QSsybHCHsZ6RlJHAlB8Xvu46ACuBzAyrVwOJpcwKtYxQmQUYievgWEDRYzIgx3o+4mhgwi3cbTdiKeABYm9JOu0GSObc1dnM0uU7pPYB0RGXBiRh5EpI7eOkZR6p4KvGAJllKw9EfezhBG95/g8Wsy4jpGEHWM/1Pcja0S8rcjIYlj3uONXN5sysjbw9XkhoHQjrI4XMJFNo3KlLkoVQPkHZ4nlk/4DaRvWirogpbVYBy0WX1lkWCuXdaNIKs7whgQsetUK9FSB18pP3Tyh2Z0pczRTYWx9ERjYpInaTKJsm7pVh2cTfaFmVThT1b50Q3TKRbSzaZ5gLYtnM0axSpBizc0YhSsyEsOxVi7zE0uKLSh7AxJFM8hdIp7DutgxTEVttEEcl5M775Q1OK5XRibTBSrZpdpXKCyVmF8evQ2fMKKUrzTfeYzdEN1qiRlReGWMhGSB05PRkwBkFucVGLF7l4qRwlZE0B6L1WK8RUORkHmtWoJclkPiYByau5FRhcqViFk1w4zi/Rw6EwKxCZEYtdhTjYxicSAz8g6jus+H8rSG+cZISCZee8oo7edgL0WMujwnC+YbGbU4/FqBDCzSbCeg66hbLqFQb5orPxH0a2wA1RjUvkKnvIy2nULpxgqdvhF4Y9ZIXbWMm5Gkms+aDK1sQq26lKzKhyEDwCPQefO1s0l0yiWuIA3qjsMAayW54TlXwmWIt4GLJZX7GulnFfq8ANXUy4c2ycKP4lquVYmVH8PCoJ1NY3l0XuNvifmpH6FEt1xCy06gcmPI6RZnIMRybDG0kZEMqiNGRhk5ZRSEDf8uC76wE+iWi6hDhXSgbAhAp1zksnWqZpRWbhl3J+lAcYFzXUi0tko3VJd4M0bSqQqQ0Gph0baTWBqd188mA2qdJ71mrVxGy6xj5EtNxUlmSkJXbelXRpYZGX0mUvI3ZyTduWvlEjFizUQqElfLBRRmApkl7yOTFCEfGBsZ8c8KyToSz9dERmJMI3/SxzJkaNkJLI8vIOMqYXkuFxzd+F51UJg2KkczKoiRhKDCKI7+k6LC6CNnKIQRa2DKSD2eoPqd1Np0y2U1YrmR1vmA1fFltO1kw6MXr84H+j5W5vWtjBfQspN6gsmpR1aXqYXo7lMcF/TvUJxPxSvi0uasulMRkhTXJFoGP8xkNo1xPVLxCwB65aqmoSQlSid2bFqLtft0C5QISj5QZkAKU6jxR0bz5/AhaGGMfI7CRNe2lU3h0vAMfKAJV+JCro4vs+gDPdmlkSwW+aSxJCKfEAu3pLEJADHhU9P5WoU3rUbk/0ZGPGUUxcyMVX2NXU0GE+Jl1qIP5KatwqR4ZJLmk/6ByMhvZGTb+mwtO4VLg1PwCByOUeixVi2jZdsa4GglIReSBc6+aYgY5CDajBFtBBEer8yIPmFhJ1AxIzEsvaqDlploaEbCSMRHKTKUXpg61Bx6y+U9fMWg4/Q5JDMFZYRNGBVmApcGZwBAGVWupPfG2hwdosnVAFpsF7WaoIy8rreUER0oCaPgkr4lmYdBBYi5bbEzENdvv6JwUUV93lPGSLu7RWZzk73v4Vu/0M0vtFtcMioRnwXVBNALYSEtyGWtsdorveBXR4kFp3EaTDwdSPwij4AmPkEhG0OpnZadULU6HV0mdQ4x7g3UeQgRi5Lx8YassSwGtnT6jwyWrfk0LWyL03RS10H1HmvVMiazGRrXXy2jlU1uyijj+nthI7/omePN68bQ1OvISG50E2FWDDRVG5LAGlQcQ6A0LHXSklptQdkIuQqPTlUq2QXAJcDxBLWIhXdSfKaGTRxcE72eJqOKOdOvzFDD4GQ+w4o+vTdhJEaTGCVl4gaNMKHJyMBxkZwP8Tb1zRk5EnsDFYyJ6Fv7EkXWRq9abmhvFacexfOo+bOUfgwZSSdzNKPQaDYwouIr6LpOGcWyAaM/d61awVQ+g9INOc0+kWhaLKbCKyNcgZFN/rsUZnnINQx+AyMpBCwsG7Rkilcd6PDuVcto58IoR+lHqitlyPUayWrNjLLjD+z/1cmtxaQsICr+KJIinjh8Q9RfcbnJ7aVTTSDHdFFs35X6dqkslHmbgb+zjEm3JsPS+AIm8xmIaKMyJdeti+cj1XI0c9Kr4SL1OnD85zi+5JumIVWOtJHTRhq5dCUdNW9Nhk65iKHrYyKbZkMUGeloNG3OAlvjyAzg8mQTZxtKT0YU9KTQJ+MXangIa4yjJRSwxmJpfAFT+aw+O5Kfm84lCbzpLJLOX66sFaMpeop0zAqrKzOKsToxsuiUl3lwzTsw0oNDnjV2mhpmFIxMr8p0yIzqMEEa3mL/h7XZpozAdQ/T+VZIOnIzRvFAXMeItQLhIR3I4pFZE/umpMFO3iXthzggKWMBv1NeRumHaryajKK+po1+xiTGgQxE1EzI85E5KpszwjswoirNlfFFTBVb9RCX9SXDqH3CyAwnx7ZXrobKj2IcLD8EFjnHUTpARawWJHNBJ1rFU6gkvrYcX2W2pV184j5ZTu2IjhGr3UAuo53EqB5ARDGKa6mLUhVvQqfVhIZd0Dhmnar4jMk0bGjbaYj4IwYqDpyhKUQiilo+mUs3wqDqoletoPLlBkaiSWhhGuIcTFmkBhalH/PX089uMGJOovHIQtL6DKARDvQ4CzNywiimp02DEaXDMuZr2FWVNLYq/5yZCghoZ9O8wCMjMqDEaOyHHMcbPSDGzGitWonpus0YhUorcpuMZLjLmL+efnbLTiaMcqqchXQos/Duo4Ymbd2NdeQGMBBX3G7KiOaFbGRU+1rZUvaOskcT2TQCYioz43UkwuPYDxGDLKvrqF91sVauNMLAkPxN2fySdo33lMTO75LXGVU5r1tHtlBjLh6+hG0bGXn06i4KO8lzVeL60RYECV/4cC+ywmR3feTGf95rX5yUhWtgVbACu/Ny85SUispJJNoEAK2UjLX9VSPtpF2C/Lu4dvI9h3WPFqil69tKN1IPQ1w6GftG/x70dBArCsQ5FbUvYZEhmHj7tZwK4lJKSpTKhanPQQaSUJn7KoyxaGdTWCuXdXKSnHwyA1LrN5LPI9WO6SBfmtMY72MQUS2KbYFj+OQineR70o3vYHXbofLjd2GE6NUhpketTRiZZI4Hu/zZekY2ZSSVrFRR2K9WYUzGjJZQ2AkV9SpP1y4gBESvdD0j8cz+nozYAxRBV4wIdUUTI+cd6lBiIptOGIXkRIZuiPTSJcBQ6hQ5aj/WzIFsNBmiLN+P2gAKSNm5ajUIjdvUWnaCxF87AekkrtwIksndnBF5WlYzVJpeaDIKQb1SyR7J/oiDmGlPDyvqHCdG5Ay0s6m4VyHeS64/Ef3WyJaD+v8v7AySG7lhKIoPkq2JnSl7MuVZJbfIFbLJKXKJnCE39cIZJ9LEstTdJH4WJMjuxFOz00LFkl4RBPAJgI+HcCun5bPYpiaiq+qbjei6hW8Ga3fMrmS7Z6nfjX3Ghacqo2Ft1GBAIMf5Sfy60esjFKHV3I8wks2QbHOf7AeRf/ZiIPVQsIePbex5yymlGVE9coby7NrJax7dmiQl6qG3t7tnHgVYQ63YMcJmQrr8lxH7bcJQq0d47sefaw/H+Ul83qenYIDWPokdI24YjXZoD6/d28x26amHbRk1j71jxL06Xxld5JJfxGeCVEZTYzTW9MNgMKqGKRtGblhbRv4/Y2ckG0bjcBGRzvg4/7lj5M9bnNcvG0bYMLINo9B/c2W0yGLXfjvnTzb+n5EMjp4OtxXnUkfh9VkuUvuZjq293Sx/gxG7bQ1GzYF0Rtajr7rPPNUackG1m+oMTvOTeLGV25qxyCX/s8kYRlmBp2Lza37EL7/9/OvDj3d/TN/Hn+b1wvubB53SpFETSinW81erj8V6MVZdEQS0uoOq4DKEgKVcGZHQPBVF6tD0qAlk7THPJVuKBz2d/yopRTUjfSOsZZEpHZDLKqVk3t1+1LWsVPcFAAoLtfVEQBV9ZkS7djUaEyZRVeSSaVLQtBKqBhhJACi29HUognmZ7WX5mwFRRAkaqO3EBiDX9cIfbj5pSulNRrHP2nRGUrt6KyMKIc6ohrIGVkigkEkTbDBiigeczs8lpUmtGFVVBBArWVKasJZFrJB3Nx90tcFIABiNvbdGAZr19KFdrTJikvAVRmyncLaVoTMC5uViL8uRAVGohOwZYV4v9uHmk6Y0adAAK7ZhZBJ0eMlq0UKFfoVRrBurqX0mxqQTjEYKUUphihNO588lpUNjFOoeaIyWvIhQ+P67e81vMmp6CgCaEVDsGSUJGt5gpGi1UTtGIsDrfC7e+k4lYCA2jJb1ave3D5piZVRKaQVDbFpBEArruJkWnqoo94wUS1nYZrh0r2l0RiTFYCwMSPjy+rxn1KKiFBOWfBWVyNt37zVb3jKS+Tw/vjyvv/8Lp1T9JBHZ0lkAAAAASUVORK5CYII="}]}
