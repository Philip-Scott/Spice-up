{"current-slide":0, "aspect-ratio":-1, "slides": [{"background-color":"linear-gradient(to bottom, #3689e6 0%, #4d158a 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/black-linen.png" , "items": [{"x": -633,"y": 439,"w": 2801,"h": 403,"type":"text","text": "","text-data":"{title}","font": "open sans","color": "#f4f4f4","font-size": 28, "font-style":"regular", "justification": 1 }, {"x": -636,"y": 750,"w": 2810,"h": 220,"type":"text","text": "","text-data": "{subtitle}","font": "open sans","color": "#64baff","font-size": 21, "font-style":"light italic", "justification": 1 }], "preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nGy9TZJsy84s5FLEyqp97tcAevAwYwL0aDIEzBgPM+ANjnFgdIF7T1XlWiHRkLsi6j622bG9T/1kroxQSC6XS2H/6X/6X/+Xz//6v/vP4/rznzCmAchct5uNzPXA5gVkJtyR6zYbL8T9DcBhDiAS5p7wgXhud/eobyRi3ebzM4FEPo/562NlLEcuZCJtXECGIRYwZsZ9u48RyDD4qPcFDBkAAPgAgMRaBgQwX5mx3ILPh0zzYXm/zcas1xkXzJDx3DBzwN2QmcgEzIFcgE8gA/G8zcesZ3MHzBHvL/MxAQBr3TDzdB+WZmn1VAbzjHWbAWnzA4hliEBapsEt4oGPKzMD5sMywsyQmZnmA4hlEQtuA5ELNq7EWm5mCQNsXpkR/LkHfn0CzwMMT/OJXI8BljDUWgKw15/Mny+DATBDZiRgMHNDBACtaX12rm+mft/Mah8tEQ8/KhC5MOZnZjwGGLi4Zj4DEQYfiVwGG8hclus2nx+BCMCAdf/YuD4y1zK4ISPSfBiQMJ/IWDDzxJhALOS6HeZp5v2MWDfgo54pE/3HAJhnPrebj8y1YHPUZwAsY8HGRLy/AXPYGMB6YD4zDYYVMLeEOfS8GLPeIxZsfmbG27ACGCMBM6C+Bx/I5zGbQ+sA2ln9jFnZbwRiPfAx6lkz3DITJvudhuen9iLTfb4iM5HrDRuvOi+ZCau1r/eeQC7a7wttVwbE/WPuox4z7oQPONzSLQ0GGCwz02JZmqeNCUTQfpHIwHp//Z8///f/9b/Nz//qv/3fP/6H//l/vO8b4/pEPG8YkucUsPkCMur/1w27/gA//4Q2L3nYbLyA+29gftQhBJA//wJef8F8IJ83wNeqxX+AcSHXXe8zJvD+Aq5PxHpgY8BsICOAfFAbf8HMEfd3+a/rA/n8IAHYuGA+EesG4oG9/oG4v+t1/UL8/L/w+VELDANQZ6sM6EJmIO8vhF8wd8gE8/7GcseYn8D9hQSwYHzdAZ56gJ8v66Ah7h/YuBAZ9ZnnR71rHYD62QiUE36AXFgRgBns+kTGw+8PuF/1/7mATOS4ev1D62kGmCPXDXMHxgdy/dS6jVn25V72Gwt02PD5gYwHMIPPF7DuekatqfF3nh86qR/k/KDBX3X4fv4F//iPeu9xIe4v2LgA7gXmJzIDZgZ73sD1CcvgcwTgExkP/PqDuL/qfVBnzTLokPj7g2uxFsbrD+J5A+51mMdVrxkPYAOG5Ne4Bxn1XO9/lWOiHdr1+csmYc59esOvP4xXtw4rHRr49dU2leuu388oZ2Tj1775uJAA7cxhfiHXuyxxXHLqyPXAX3/Vz41X2fz7XxivP8igZVrFAQag+r33F2K+2unCDPn8YMFqn+8vmA+sDPh4IZ3PuN7IjPoZBo64v+HXH+Tzg9ec/w3wf/znCRv//f39hczEAp31uvfGw2lY9ZDr5+/+N8AADa9DCqcjLcNEgh++DDS44ZmrNn/Uz9fXAPgF2AQsAAyYX4jnb5hPwBhEzHrTzF9Iz3JETgfuFxJexjJeO+iMD8AGjTDKUZgjLWE26sWFNmzy4wV/x/itMtQKFBOAIVbQuTgM1huViYpOFQ7LYPk6GQkE6nMJ5GAAXq8BeP1nVu8zXrWJmXWoXh+I5wfmtUZy2mYTaYlChPwcbrUWVvtl8wNYDzIeHkQv52mj1nMFnecDs1mOZj31DOBr2ixQVt5qOyCj0cLrWVGHPBmlM/n/ayHWXdZmhlwPMhOxFnItLCMKzKyDho0AM959kDNWHdyK4rCo/crnQcQ3bH7C8t4HOhNrfZeNHnsTEUDo0LVpA0kQuu56lgLM/DxGJxztuMtO6zXcefjXu/YlF5Lny8YH3/oqMPj80KaciKfsF361jZRdDyRofyjUk8+7bOD5QSHHUevltu2XAB1eNisHXXuUtDf9bYqlyCjbXBiYr8//NMvgGMH1JwI2XuXJzZCRvSGwMhCzMjBw03xe9EpZH5oLWge4FsHHRKUDA4nFnz2iPL2aEfZhXCBMr7/1utwYGVTBsYcH3SoaxsPXLq9tsfi5BgjV6nvwcjzmFUWYQvn8qEPnTx3KcVV0eL3q8JjBvQ5n/XvBjIfdZ0Vdp9Nx344hHiTXXJFnmHMPF51CdPTw+arftwEM59ouvv5oJ6LP5D4KjYwX1nrX+8gA4DR8OkLUZ1jxwHgoCn2A+5G9Fwar/Vu3LAlIA7xew+CIuGE+4fx8kUlH5fWclr3nzmc3n9vxWSFMH69GO2azobvQIzJg85N2TUSFVeup9Zgf/MxoO6gDlLTfsQ9zgiluBQwzI7JMrq2cglXA8x1c6rXx6/+1h2azn8nG5Fla7VzcBxYPOejQzCciFoxrDqJYI2Jyn7VHkdyTi+djVhZgXufWC7W70859wjNh80I+P2WrY9Q54D7VuaLjG6/63O5lg/MTM9djxUHQnaCgi42JtMqxMgMWC/G8CVUfBGJHZAsiiAWbhoh3vda66yHMkc+N5GHPDCD4vVx87wWsBRvBiLUKMTw396JgakWqh85jyFfDjIeCr+8+Nxx+blhWVC3oK4e39xnxcNFRXnctGlbQ4YGf46FDw974pFfuqMT30EZEANP3/6/7WO/Yz4SEWx1Wh+tL5eT4OZU21SEcRHU/ALz8OJ8pn3cBNIahpJEb0R54+PJ5A4tQP990vLlhtzGFzEREIO6vcm4KGKvSKu0tMolELmC9Ee+/uRb13JaJfO6KpgDgD7AeYGTZ23MXenkKGmfSMZoj7x9gBOL9Rf5p8JD5r8gd9zc8XzzUYPQsx+DzVZ/HGGljEdrTgbgz0usQPbSHu38un5sIIDvl6PTEr3I+q9LIfO6KmWvBr8+K1kE0EEGHgNpLofKsT1KUwPE1pYzBTyoYRPu1SJhxX0L2SyeUs57zucvJt10LTfB9FCRQZwQZPINpc4yZ9vpHRfzxqh96GSERPRtkyAM+PxH2VdFtfu6DCwCoyFL56oNUygCD+YCPDwTeACraVOQdjNR+cAU8/OZIK14AuZiX7hQhM3gI5o7UXMSUt7TBgyivzjwzFl/bNyxbD9/7WDwzGsLDFETE6M4dyz+8Yf5n/0wGkGP/TH8tG3I2RC/2iQYP+PUXXycqOhA1JNGTYD3kVJuU9HYqG0/zz6KT8+tY78m9KTRo81VcixOh+SC6+UTn+0z/kD+VciFg+SpnNbRXIEz/gM9AEcRXpbWMguPFiGsD6fX8Pq5KCWCw+dFGXz+H3mf/nJ1+xCqbEwFoSODjPzpKoyN5Asrnc3/eIoSNadygE5BDQae8MIeT08NQymGVytXCHmtugE0+c6EsMNUSwiwTloOhYyMPIgdgRkTLZ5TtFHIpx9QRxRwAg47IYP1/BtJWozW9VlqWY4Mh7x9yZcGzFsCgUzGi6n5hQ2/M9lj6e0OvzGdvAKOxYFQZbe5c9DBqI4m1F6p+toyYORUEs2N7PDqFZsNFvBLVFGGr1+WBFFyTI+CBF3ln5CGA3J83F8nGuz3sji6Dac/YEBQ68A8N9drrQidpY+yNa2JstIMBCora8fquQ6LnJpLqzxzRTiHlAARjUdEIjMidzlQSjU4j6bySKUUfplgAotNB/X4Rx28a9tz7JccQTztz7VelXHc7KHCt+g8RSKVe/D1VaXIh18+OjhntG+vnZUMPRFfXhydXJHvR5+Bn3O9FuxZ3Q4RS/EjudZJNWQWvIqKz38vE1eiP0X4RDDjea1L2zMBg6OerCP7w31bnQY6594A833rTDooCkNPAcWbzWLNO0c3ptCbPTbTdKAjKcRqdrI1XB2AhRkcE4v4pyMEPVy9AT8TFyPX0AUo9DA+GKhrOvP5cUKxa1Fqwi9GaqQkjnPuE284ZxTv4qEhgWQanhzd4H1YbryKTROIwh5VB1utclT8OemJFFjqU+m82z9JopVMLetgg2aYDZl7pCqs2Yt7lSHOtXoPaMFZ/SKiBxtaHns9XRgDuCY9C7DVP/m4bnI8iLpmbmg+M+afz+/55v/ozFTFqB5fCiM71NT4vRKqOj+Jo1k1DRBuuEXHqPSB+SKkhjgNMlImkvQCkMpLBRzn2i5+d0ZRocB/yBZGNnTb0utfa9+FOVIrcAUBoYABp5WCxbYBcMN/z+KwiG8V30PmfNtmfW4eTn9X8VTYI589yrVntaOTgRVCKQzQ4bFxwv7gf0euugCg7zlidnphfx+vWOpV97/eWXXeqoyoKnYgcV/FNnjOyyJQEgFvR7NlRZOxcPNZdHBG5iIzvPrTwiVg/MCtoWgGniKvMefwOS4eqO+dCrAXYjbx/EGTVY93A86amAwX3FG3bkxe/0nCW8CnEXseCxYN43kwTJnx+1GsSQpZDrBJlrrtSq/XG+qkoUN+/EfLAXmsTsGag8fwg101Cz6r6s6TrGIyA2Qc840Hcgo719XgeiAj08WI1ajYCkEPJdQPXJ/NwIja+V6JKnGmGRQeeq6JlZhTEF2qhUaWcfaKqQ1F8SvFTH3ud11PPEauCCwA8Va3IWMifiqbr/cXNyapsvP8WiKtSOfcDsRDckyKjnTl9EE3dVf0Q6RoJ4Gkiu6LhxxHZA3nvfD3jC3Z9MIgI7RQpW2vp20lTp5BPcM1UcXkYK7zRrSKxz08IjYn0zeeNGA9Kc/QGcmG9q1xpKhNrz2G0uXelJ7GQtO1yfoVEl/ZJZVyzkgT4RFoU2pCTIVcUzw+Mr5vPD22MlaOo9eYnLcew3uVABqsz66s+CwONuyOfH3MnnGwvqHSApR8wr6qS17sjc8Md1rBT/7btgTvaJ6spShPMjsga/bNdxuFClaGMzVNw4zoiP2L29fViottT0ou6X/SkREjKL2OV5z7Y7Xi+O+WRMXVeSFRlJFYb6vJzllPgyWgug5FYh52R71c1RwbBQ9zIbj18Br5Wk2na/2d/HjAdMaeDYErFPNhb/1LoK9bNj6VKgXNPRbipjAuc3M1eVzpjpkDiYKx1I7VmZjvYKPXo/YFek1B7PeXsVNmiE8m1+P756z99/YyuQpbFNaCdGbIOczNwTJF26iRtESsJqZRBKFawH9zrOPbsQNPtrGpvqnpxaQH6c+j7WhcQgZz2YGboigfT7raHjEZa4pLK0bwbGW0+RtmA0hLb+0JE2Wtx/iHak/ZjgmXLMjVHCfxibwKFLpmBMT8L/hA6FSH2zbKQI8erUwwfAOYHfHyUV8socdFE544mZ2JF7vTB5eaa9AUiF1HQi0W/IsSenzY6pSWJd0dp08Y8b9h8Ve4o/mBIo0DdRUY9rw4eUCW7AyaqLu46UEYhlBYXciIPIyrThCM69fOOa1ebTrGYyl/JUmindQGqFyDY3YeIOXalbAfRyc+Xz3s/mznTPtvvmyAKpBiMz2SwJo1LZPZD5PMmj+mHww24zSp5i1cxb1GZDH/rCV6FBm22Tfl4gSrYKnUCSI99eERqkviOLuMLXntXhMzrubqCNj/qPbzIVhtVMXP/rZeAOcZ4Ia3sQVyL+4UciVjZtisHDUSdpK7woT5frI7q5Yis1+20X5N2QyrWI+XLVXxblcSvrk4Vf0RBGtNXtxckpENmVb3OfYxA3m/AZq9pa1UiYMMq6NK5dXDwSdVOBuK5MV5/tacv5d+r8+vamFWbCVYU7h8eICrBQOZay9gwcmwvFtwAenBTWsNc1m0g8MD9tVEErHPiJpF08EQoEtLJ6QBWB2eQUR4X34/OjIc2hXaAJuJAZaXZwJD6EJVqWQKuPJXCnJAxjmtvQOpg0su7oQS2PFjtyY/3Fxklxz0udBnLBiki68guTgKWLUCLVBrAXfALZtFwvXkRPOSYNokJVmV8vpCMiFJ9RnwfqKIcvs+P2uOnEKdhIyWV4Bii0JoTWO+jbEdrYHZh82FGSPzmS0Sx9XyGODQkyTL7eP2BOIkSQ4ndZ1BSaZP6CuTqwy5EKHWm2QTsKdWyEOQqTqVtgmtWlZPiKZw6CbdJdFklXb/+QGnILpfy36OCSTzvsquUmxevURUsZ2UR49VBBRRO1RpfO6glSmFMVeZGz+KKSjcDM1g8QFrpLk4Owybg2bzGRESWlxMMjS5Rlkf+6YNcXnq1BxchKu8Xz0/pMAz1u88b/voHjWGr6IpnSNhQvixyiocOVTfvfJ2HVSpFleY2B7CAFPQMHrBSaIIGLHKxnQtsS5LJEMsb75IVS6mMzj5ejEY/teDcAJ8fiGWdx6oHocjZMl6ffyrCUwHq44NwMEpjQKhXG55EPfUsPksIFg0ljwMmh8HzUAbBspqNqvPLWXc+sFO/cp7ZHEkpNsn5mFdU44HvqlOnHUfZlihCRrxT16dFbO1YWDnqaM7opgierJAlRKgLYt/NGyjwKcU1EeaKhj72/3O/xR/pEIKOxjJoZ0yXDaULyrUJ4EZ/KB3H/CBC/U06K01QyhLik/gsotyakNQzUSzIb9aKqnydpRvK501eAQyaA4ngURD6YpDyUfY7Zzs5n58wdz7/i7+fDMzW6UxmwsdHrZET3c5XzMhl9pDgIByL5w1bD9OLsTdrFbyP+wuwUQqviCLJVC2IQimSdIsUq8X+KdhFgxSBIuPO9a7i0pLoperk8byRg2RUV2kCeAHxsCmIhF6doQc2mOpQMptR0S/k4NwBplBi1uN5wzOBAeD+QcTDFKh085Fv5Jsoqyny0WRdn0XsnFSa+/X+V38/40GICDTrQ2hjYv38Ez5fzfBrA+P5gRhyz0A1p716fVX3P2XhRQ4n4tmqxJNoWz//gs3XRnYRRYjxAKta3+U1nyTuchs6D1r9XCkV4/3F9PXuzyZNQT5vhMjolFT8YYoDlBiMeg4jUQjUPj1vkoCFAqpHKGCLB4ypSBGAp9w/AUqukcHUmSgSoEjsDfFB+bybN8lV5DYTRCIdx7q/6Js3FyCHftpvPnc1BxJZbQRcZfJ4ShBpJKIB671vtS3A31HJvLQ3EV8dsJLnBBD98ex9WXe91/vvDhhdPCVKQyZclQ85ZpGi8wN5f9tsyO6zo1TBSwmtrOGe++xcU94RDh5IBmJGbMuJtIqUqjDYuDDak5L3GAMS7CCjjFfSU3OkD4yPo7wkchSJ8fEPLNgmxDKAMWF4Ybz+Ktbe2Cy1invxcW2t1ARhrSAj4ThJWlc+SvWljU/uHKOV6bNMODkIZ84ZLD+qUtMpDiG2okhHhFlIYrwmn7MgpyoS5lmNluIpFmvnNoG5U5h4fwHum3vhM2QslpipeFxv2PWnHI5Npl3FO3V0Fqej6ti40OU+PxrTjBJ6L0P0+eJ+qq9BknMHrnKKhgsSUslBST9QPFds+NxoYfbzgNU0E/AhB4AMYH7u6Crob14nxCdMnJy4inFR/0qCnYjUnBzKoAZhfGC0PJ2Hv99+IkAnKUm6DeTcqbKcE7xQqc9K6SMeBuWqsti4MK4/R//PRPpF8x/1bx9wY+PnnE0VdJsGgGSKl3zWcb3aAeLk0bq8e5UMn8HTxwuBd50ZnzkNSLHAse4SLskfy9AVSRPwSTJz3Y0oZEz6I8gVj8iwhVgPhl/0zKwczFfDT89s4lDerA1DrLQWO6scsH7+iRC8622rSLXef0N9JAmWvHJhSalH02gHEkdfBpudoPQJ2Ko+CLm8IHl09z7cP4hB61UHYwbieVpTUHmpIXH/Sifi/mpiyiSgApGTIlc6cn1XV2aT5ovEp5xYOaRY79axNLzvvgamBu4la8gHwATANMkG4vnCwF9tTBsyr5ZiG3tQqqy8EagiXYuu1qkcDHIR1TwV93d9TX0bTHMynv5MSgFUYgVZHTNHQO0Cue1X+oyHUmcDIh8U8evY/RtrP6e4NdvpVtwq7VJYFfN3WZ7cVOYDW1USdp0bppF1MGW71ntmubCICtu+U2tX9pu5YDHY2U6xoBxPHgpmOQBVyI7KFY0R5kSr5qQLPst2fFDbku2cyiQXMGovorhJn7CaiQBWKzr/QkXcKltSk9CcwTdaQSmiqnOqAfMtn1WlQQ1jgtuqDzdr37l4RUOL1YvSEeV5U3sgp1BkasYCJvskqKnw1z/osZ0QrbQBFbHpFCgTrj4X5dPseWHuvZ43VGZK9rEUDyDZuQ7sAoaUgPFbF2EDHQIzEesNn1b2Ic1JRHU1xkJCZbTVcFm18NMZ5/10tUrEY9z/gnQDiECAwhoRl5RH16FMwMqJiuMp3mQbYI0X+Gn421wH90maBHQlZiDASpcUnuSYqlLxAMl8+bARyA6alOW+1UCAIkLp5F32AxLWLL0aka94Nbg1QrY8SWFyNYm247Y9BoZ4tqMoInwHo+bqRiG1U1kr7s2OcmV3nTKVs8jS9mHbr6QLcZfGwT/+oz6HU2X5/NT7DOO+JW3xu51DdV9vesB8VLrEfejuW1Zoal1QewKDj9F7CephYt3VT52RM9ftUJ5KKNMEVwYchN4sd2Z7sWxyplDAKjhJj1qVDypAhUTkXNbd3YzJhy7PXaWboCDHxwe882MnaXgd8GwgFkuyRBtuA5h/iIgWIbDKkYwqoeaarNQqATXgiAnWwBsn4SiHZj4KygLbeCrX4XsC1Y0p6L3l3VV2nmzPZteqnI3IWNeh2j0hznkUu5tRbAKZa9slUGcFpVO18So0x9k4LftGNa3ZmIhHRg1+H1UVeX3uPD5u+JhYTzUJNlmsAyajk6NkCtBNTchCD+SxkCKzQQckR7QQ73/y8Hu3AySb4OqAPG3UW0LugNN+1aRmu3LQmpCk3kIcTzywy3bvxlVCLwn2KlUhAmlC/dmHTvwXA1CpUZn2zQ/yck+nPdWNS6WlyqzdL6KZF5Qt2JZbV3WFeye6zHfJWvYlB+1efVLqStWf7uJW2qVg7keflKFSN1jZiBPHZXmFhubRqjb2KST6wHe/e8uHWV6jVLYIL+Z93KCWy0ZCCs4Nl1Fed0nYFQDnQpwyVIl8NDdBkXtD3WJ7RQCGhD0t1d1GmmxPFvkIMuKpMl4sRlFJ3hU19xrVm9TnlEwaEew9YVrWwiT0hvTPMQ2L91f/bFLVqG5X68+9P2tHaX2ty4RcH1YfSs/wAiJJxHkb+Wblx4bUkqAn+jk1eEgEKjJJbgJu6jGgEwbwa64DrPfW5FDzdx+FZPxCCyo9lqXqeck3dE8DHQtL9eXA+V4k+oLqTNmm0hqDfh4MhJRE+4RBpXDfDiH/zX7lqPJYp6zPoWrDThfVoAWoTSA7xagUV/L1YEDtpkKKH/V9BYOuFvXrPjwj/vsZdQYkdadt914d56HXA5oz8ub7P9uuaesJ5GzNuUggHyVEYg3ZfGCMf2A9X3wgzhWQp9y7D9WwDShk4BfUx+/zdRBd6Lbo/h6so7iRzOlauks3Ufm8m/9agEptVHPns8eG/fV4ju449AGL0dFXJc7+HqOJcuMyoP1+/95opQhn6o/oDVYrOjrflgfv9zlk4eIEMiXLVlnQdnooQpQIoZ6N6IL2spFHlWi3jmVrJBo2o0q+Kr/V4JwXpOSU+4gI+CQRrPfTftvR9av2fKDhb5NuPlsvkLnIvVTru9GnmF+N6iy9kGxHTonjYu+VpoBZoTKHdSeq1sTmP5obQXJWy5iF8jJQOf1ukFOkRV7kOQopVrRtoX2nVjhJYTDVNVS6ymlwvZqtk8G23zjmwSjYKjiIjzOvWRQSbIWcb9Lhys6pZLVDX3LwF4XuiGZghWz0/UFyH47MG8izgzrOIQx14CGZd0rHrtIKD5xJpixiLwm5wQ+x8892Dpz81F2bmgSVVaLZpTdqLA5UkCEOoV6zSJoNvXrBFNEz9oIq6kYZVxlM7t4GHEScyk9LvQuK3oK7qqPf++efm6Xi0qKIRN2qQXEXREiounuo10NRIJ563/v7+NzMSaVToHPMM88+OJ9GWILmcixMDZDrQAlo44LKsop25o3SjDUCSIDWqk9vx6z1FlIz7MbCstVN3O33ZQ6tkQCjmvy2ZoQ/S/7B1ZGrKpwPHlQhER28wUYsWUtxCCKm+8C37kQO+erf0JgAOfRdHaFAiqrJ7kHRXp6clpCaELKNw97fe/9q8xt1CUkCCY16jOdu5xjv79obtTmQt5NkoV7j3Xxgj2ZkugHwvBFtqER8lr438o1fNpGx4DggKzLZaVYG8u8daeojUOTs6KTuyFiUESsvJswJ1YxpBISjmvZkSk9+QeXNH/RB/SXasYKPSiM6ZdAB0KYINtJZ8TXbwOh5z/y7vrU98z4oQENcq8YnmBMREXbb/P0zkyXiHnYyKHneKZnB4Uz7hPCMBxnkIsrxvTfncsJIHcb+GvfMJuEona4OnRh+lcj6+Y80K9linoAdnE07h3MNfacl5aiv3gfgcGghgjyPPDrbMXdKq45YlVH5Ci1w0usIGemwR1Ya17ajNLQ+m9EO6jPx5+201eyUBJFtKw3LM+t3SKDWcCBJyqvPSD8rla3WDFnNcWWvRHo2e80kbtQ+/rLfY2SjnlNrvwlk8g1yxPwemazDQdE5u0rglEwAlEaMthG1T8hJziqNfHPSkaK0yojN1wIpgc3VhpvXP5osSlTpygiLY+nnaRDAcaDr79AeHZLwbsaKVV11sX5/0PJv/QzgYmhMW5s2S0ypUW6wQk00nOZWjKRosBrEur4Gp0Rko52Wc6vVHbtgq4Mmwq429+qKTP0MN1I/b+g8vvJnDpVBVSaKmf+o9VtRw5K5HiljEfwdE0hWLliqy3xI/kY/F1Q2BIBujqruUafct0hWGR0PdUT3aFTkXDzqmqBGWTGdWala7yqb27srbbGqPI6z3Jd10Nb7n/VWdwnWchnXSOlDQfpEoMq9RHqC4sZydCymF8AeNqMSbCkbA7Xv2Q11/KymYb1SLjMymyNdytRzBgs69UoAIJn5y7F1f4+0QoXEa8IZ2gl0NYXIjbBuBzOX0hjbRgyQOO53sMk+T+W3g+R3yeqRuUcqMvh3Ondog/L5rrWFYWaEQ8N2jUq6+2vnPoI6Yo4xdmegqxKph+MAACAASURBVOZMsiWDk4MEU4PvM379jLy0q5TGqNcHIUs+vjsHOQdTRpuHqOaoe/f3MpBZrL2G0jTqoKNxOrgaASftyBsIcgFGTQUnNpt5sexZBKpffwritwIzGh2ZD+T93W3vPQ6NGxHvv2EfUr3Wa0QGbN1QKz2MvTgZtX5U8OW64VQLmtXAYalcpQ5UKc3o8JMiojYGFJqI+4u9AzS4xRkGRqczqwnQjP0OjHp+zWqBj4O3iuqwLATxbihuTe6iSbmSXCabo+rvlGaDrdilFlZ7AcuQ0s0c6sr9p6oS5letL4e3VLtCxyvAdwsB7PpFJNch5XozV7ex+y26JCri1diCIGQSW5MCWIn5RD6qmqPUcFxwzi3tEnIsmK1aD/EVajaMG1hyTnT+dFwSSaq8no0y9MGLElDre6w3xvXXIUW/mdYtSvZp47kVvfn8YJp7dAusHsQnxvUXVH+3yYYZcwqY3rDxB2eHXB1cg3riEwbM3BEHYKnwSGF8lDFdnxzSGk2ICn6bVIuokmr9DqOj2X59n8h8s8NRsxGeTnMC7wMVlBH0iDQbu+TISoFG/GfnrkBN5Ga+KuIRVg04qXZpknPsalTXqHpBMhbG6y864+h7KSTk0fuVYpKk8ZglgMtoTT/oSCVWgohGRSafbTRnH0APWj6eYzdvAbBXNUONxcNf80kGU64xPxqWOlFPqRw3glGDWY1Q3IOL63euHeFGSB3IVG1X1HqATEdnwfBEBr/eufi2l9KmvDDYuLVVoDo4DrMa5qPSfw9tqoesNVSzFQc3w9h1mgs+Ej2EeaHTkXi+ywmLxGS/hT6/BhoXWM/qB7HXgT4W1yg5b3bb7yK6ELFtfiHwU+/B9VMLQqMpIlcVAcr5fPZ6qalSCKkbMwFgJJWtgFIuF8PcRKVXpyWYM5Zn3YRmvejELrFZT6oSJ1DzL71JF2v4Zf26fUAIG5uoTEDXChg1EHt8HDech1v5Wi+GUE5DyU3mnHkcWBbsSVySoJ88he/5Hls0BJJrA7q4ZeemTCVkJD6YHrH9ulMg7yi1N4q8xNHfcpJ3lQaRp1Du3NBaOTE2z/JrXbdYyA4+Q0irpkMtRktyD0f/xY560chNjXoQQcwDWwf8tSPrwQkhVu8nWAZ1r9mdTbgxpfLxIpl5zFUBGhp3FIbIcxBWl/x98N4RBbFdHfK9h9qLPjRMD0zdsuKJFAR2dQjkNDqtO8ucQquavAXZM3aKetovlPKpfyb6NQsJaEYL0BwMba6bvcj1ITcpLR5JRDS4VtsJS65ubUu/79XZhK6PF9wHZkYYCHUtDZpgjPw9r1B9ECpZptSFiZ76raaYXkCUZ6t5NruxSh+8VY4iVlE/Z8wlW8yjjZNoLN8s/ShnxUGEiUCqg1C/g32AavfqeWQcLLV1rwcANT6VoSdIBaN1FA25t6gMqbIayshG3afiXnMgzl4RdM3bEfGz0dN6CpofTiVNxG1pHcbrQpLIK3myZNxVt69ouJuQYj0wsLFuvFDderlJNO4vjuoPQPk/ozW4XvXZ6SCWehqq0rTLiOi29XhuOKrHIu6fYuDHtd+nhXB0RhEA3v2ZxFnFehOpYKe4REhQ30UvPonYVKomiTQARCNIpTY9xS0rBWvki53ygOn1Jit349d22sn08N/tF+Q6EjDalNfdLHpWHyQxzWpqmsY+8DyUkbP0LY2NeL5OI2avFzhDRjzhlhborpVJR8R9SOxyLZ07WDHB5cjnTofxGrNi3QpOYv/ZDKzk3tbQp5lmRmDpE3oIrXGIizwVeYezbi7m3+cLIl0ESXHcDCaPDHO2Bwuqao5mPYe8pvvpOdex4SBMv7qvH21M+TuKmKKT4Bqjm55HFY++DEbPGntNzlIdoyb6PeqwqN25h6S2fqX2oyLtBb8+qYkY/Zzums/ItXE1FZ1S+zoAPbRIpcdDTwJVXrT2fFYhp9ZSSCdiGjRMDkSvbUVC99ow7ajPDGp0Jl+Pc05dJUnb+8fPvVFA3cw2mM4NNTuao/tjbbP+J8IrjynENfaaANBAndY/JNOvc/8atnsffHFmMhQJwFzak0H7FcrmOXFXCTjbbhqxE8XvCsVGePUZJFJjxPfZz93EJORU9jl1qarPShtKNl/9PUoNs9+re3DUbmAwP5n6lnEnimA6YZugS26I0+dYdfZYNRgkDjhvx61K9JZOuK5cT7B0P8se4rsN1mh8ExpLp2epZziEJ3YIebygq8abnWUhzZfYEFMoXumTkIb/gv+CcCqhsdOnjQLaDqtcTzlplxS7ni0IjWONeis3WpGeYfE6wGbWs9/nTKF04E8H4rwDpHNXktA+PrcDqWPUTliCMTkbVXjcX/21PYpOLeFKM+PXPvxaN+o+xCn0FZaN1DZ5faY0Wgdk9dcoigqtts4kgyP0VFrdojGQtyo1Y63fVsgWtG9bojMu8l1cFlMIG9AlQg39D8cqlavPjw6WciobLeT+G7alCAwspnWVUyEf2Grp2KT6Tou8Bxpb2xAaESnIgXYue2lKQAFPjoV0gvvMWTr4RGaRPmBZyCWQae299ff2EJl9OHXeujSq+Y+5mPcBmRrSyoYr9hkI9oiM2Tp85fIP+vakVjEW0qm6d0BXyQl+VQPUXQSiHAFLtJK0QyXS4xkKO6/2xqqLVxRUisV7PkERz1Ot8Fqflkrn3Z+hytEcQiuoyAY2GT5M3ExNHVND23Yu0ppwDVQ2JQehpj/A2K1aOWwiaewubhzRw4V+NgeRx3uwjVnOBbGqBV2/w33Mw9BTkDsfOkDpRQj7aYk9RCezkQnYT1I/vxA3bYPIcOfsO02Ss5GT8cE1he3OywDSaC/YvNYmdtHPkEyvi4PYfSE4qoEVRPne2M+YbT9MmXPfV9Kdoedemjp8GYh0YdFRWevJb5zqnSGx1gNNGCv9SCKhSmB2fxEgrk5TyCk7eB6M13klJpvlujLJQMphv+mOiMdcRu/NmOKXutCwIbS81IkAqpyEnftFHWCnhFq5jzyf+0XDJYSC0RPepXeQ1h+CjbYjYeIwmqzmmvJ6PJCEdpmwrKYtpQlgz4Rew0VSdYnv8OYQWiqtSL03HaM+gxyO8rwlCfWeZVCvJYkyexEgH3r3ZxcUPMVNrQFQdAftMpRfPhulZG4nyyYtIwcFZDXo0RjU62ONIuY2FH5+Vwr56/VHrXcjy9lfa5gu8k1rrT4foYoox+Z2iOOW8nNvp9q2pb1mEGnbAaqKRpQKgPYrO3x+j6brtVP6e6QqIjO1dozIIn4bUfJ33fdgnlayPm/yN9rr055UvRi0ITpJEE1qeHP/3OxnM5+7gSxW4RfZqPiaQ+zYVyrILlVa1VoDdS5U0j/mdwavcSzEslENYPU7CUzESnlV5L03LtVs9EPWOpGSviZH6I3DU6sMk6qFr1bliUVHBDRtaxOJJD0T/Hl+LephK/ItRH7TCD6KKMq74piIOkaBdX91FaYMY2Ktf0GqORFTpR249yL6hEbTV42Ua37/oO47ne3J1/13jdBjWpAsyziNO0IIwbAWBUtCTcmauTnOUfj6ebrrXkdk4FlPHyKYU+eykLhZjq7BLB2RMmHG9mLdG0p4Lg3H3qdn6w4SR/RdhwiIhywrLYv7u8qEgzM41++5DwVv96yIatGunwm+tshyff4OSnQyiZpjWddK7Ma5Sgk0vUx2RGLeDmSXq543pUNg0xVKrBbx7sPXU6iICM0ACRMrw9wtBXsm6A0kiUy9TgpBHy0H8UYiEe8imJ0pQTy8MxY1DzS4P3F/QxPjypaS/mc1b6IRj30FpPQ+2m/NXUF9tgS5SJ7T9f4n/PqE2cNmwiAvcfezA6WR0Qi+XG+bsR4ztajDYXNuIQZfXC+YuYfa0HJ7UXTw6r7TVy3SWfEI5oURwBDLfcpQ0a/VOS8PB3LVs7H6IoKv4R9IAskzWnZOp7r22fFYP7pz6ibRBKfFLOfqMnJ99oMPkJLURzW2qZ6taEoi2I1X/4lDEAQ/dBpyTNW+zgtv/IXgnZhmRkX9zul/RXJWaPThOiopV9XPu9qQ2bzls/dHa9eRFkQ3Z50+E311AHP6sx+iB/eUl26nk0qHiJQSnLFqkkffreYF0KrM7DTDqQ7+zeHE/QX19Ih3Mb8Q65v2WwesUjJAYr6632b0a9n4s8VwtM9gRI6HClFxK/rcrHaJp+rnmBMW5CcgPmvzMLU0W8/QClmlXLb7r2pOLXU4GkdA4NCptqprfIWeggVpbP6g5eQkpPuyKWhMgvQ36gXKtuMe0G0jZ41A++hDAGDfYWq+J1atG8iSVWPwaInt9guZRCOMZHWYZg9ncS9GX3ddtvYgF3S1vHQP8vQqFxk7Y+P5ho2xo6wiZdY1Ba36a60AI7YdU7rH0ZFqxtF/W/jScygATmrWaxzMfIzexOYEEjzkY0duIS11zaqBTmSnIoWpXZ7wl1WF4X+VUbljcPRfrDd8fLRzLon6dRjKxX15sWNzdU7ah5idu0opdunY2ng33CYBbYzYttCXIDHlSh4EQ6I0MHm87u6yBdTh6jDjnAXZvxwZA4S33Lzyf9e1EgYgLtS8j0JTQmjKydt+h6a5E7XyQLbQyGfZpU2E7+pWfTamkRzqbLJXCqXqM19AqnxMVbENJDQZDHVAh7fDE1qrALT7aMb8g/V8Y4wPOk7nmjuDzpaAn0rc7rIGmrtTKqQJcDAHusKizmpVSAYQN5EaUfVgydZfyPhmOuSY8pjGBS60RRLHHFg3oqNLIJbINQCsFqS8NAKIyrGDJNfJcaiTsi/ySc4fSCkwSURJumxj52Q09h4oS04innelKXBk3EjsawWKdFswfNShaVIQR/SjToSKSKynGJL5wW7b2O99RFEbn50yaEMbvsvzMwqhI67y44AZG7VMfSpAhgauvqBKTXn7ecBFdt4it1xX5U86UDCKK+WrvSEygCKjVJ86OmhIX6mOoDnqOTMBZyetH52s4qp0xws0A2MTsI0wpFsZbBlIdQdnTUZzRcyro92uVu0UUk1XRTBunYzQVcTdkfWXPqdTLHJhTWgeQ3uk2YhnB44WyCXPgLQM0mjUMwfTS62jhhYjk0Q7+5kygcG0h+R2TXi7scgN6jzEw76afGr7nKMKlC5ntlMGKAijc44+O5suEJpr++0gBZzoFCRbizKowDfjeZvFQj7ftRyJyvM4Ol9TfJRWNGex3nCSQpUwVO7lsx5CfQ/J/DFzYQBQiSp4C3e9Vm12TddWOdNRt0CfJbPoA1cOibMm4yYvUHlt8SmU5noNAF5P3fy+b8UuI5CgJdeNeL5Rk6kupk339sxAR454frBsV1+0JjZIxvGeh0BC8mM8O13KeNjAQ38qqE60Emzeiee7I3GncWYH8jOs+++GxsWR/FR04vtF/r61LJGbxwB4ZeGi46to57GKq5p/sDSctluXuee6NhISCu0cfN1flFvXwVSe72ys69fJAPLmTMgPfp2DZHi4pRgFuQiAZNy4gBVs1LNuPqOnBob1fR5gRWJXY3SVX7REIMk9lQZibZtjEEIm51YmgxK6sS3yjTGzHUES/TUfgkP8pHSDB1jXYnoH68R6/6vteVx/EJkdIMTNdel6vYlGsa/l1FRzNbjRRqUNKftVpWZzYaZqns86C158ll8fyPvL5hgvYEzaG3UMwdyVfRDVuvqBeL7oOYGhfgAALTlVnovE8KsUkj7gdtEIVsFfd8Sq+woybrhH5f0cNKK6eB9qnzQ03USlaJpwWE07pnLODPDLN3HGQT2Dg2k0qk4RtiB8sh9CE8A1iu3q6LcHuUgjorkG7KRsmMfoOOoOkYh7t1Azmm0iVWXWcnI+P7Duvwnbr7rhzTVXcg9s7TSk8rSK8OVC+RkrrVv3F3z8AcZGVLlhBFRhSM5nqCjLVmUUYz/8BZ8feH7+H5i9mCq+gHGTVF00ldkOQJcwxfqu/YammVcyVE182NB9oo0ZskGiLW/kpdycowNVRXKiroOTaYTkSiXohOnQsj4YhYBVKjQ79gjWl1y5DWBs5abTXkC7T5vFkZF/q8/3aiS+BXTkQZQysJTrNqokvZ6qLPmAvf5RgcxGOx2bnxUoWkhXaCAOzZM6jM/p6LJzIaROBzmQCFBquy9ezgz4q74f467RjPMzZ8Rj4L0hxZqql95qmpQrB6M+gTCpJg/rb977EQ+WZk8w6noG0ipfG9efeg0DPTIYKR4g/66Hpqgr840tXgnEQHlpGpo2tSOzRXvckp8fAh8aFzKPlnvwsNXpiXhDV/fFEal3TZzy4KV7Oi4e0iLC1vODMa2DW3EKu41bN4sVQ31M0IL0ImyrjgU4GfL1BvBuhWdEqQtXfm0ojWM6mFqolQZEIOMHv3pbVN4DugcHfC691iLMt1mvt+4vSJi2ni/4XFj3N6ZXM16nr+vZBCdLkMUzvUoxP0qmHvjpyN2SZqWN5EDK6eaRjknQpKna0UOdNZpfYr3g3I/taPlz6918V4TmfDx1r0pzTwHJywEAukxIiFOXJmfAWA3UJHUR4ruNnX4BBjN+bRw9UfUhkWshXeMYnLZUr1PtAvvCpBhKJ9feM0rIxa9l/tT3FOAonkswpYtV3bexg0jcP/DrqGbm0w47rJDYNFioAQjKvX0z6vq4AHUNun+SG4hAR/vqkLygkeywGqahiFjvw755B3TXpeervDyYr/MdNQoP5AVWPJ3PS+RigZrO7YMVTzsikO7OGBiT9z2Y5lUU01+RX95+O4lTZ9+lPL8ABA81iUuOn/MefCNjIIyORV1BIbV8CBu5iaA8OiDR1FbR+VDHLstlzS8MdM5oIuYUXbZSNVQ50ZUyXX1xJEviYub33I3q2FXfSInD5n4fr7UWx1NEaiGJcVV0XqHIlx39C+kxarGapFJuZKLl0pLgg/9msAF5qG6/bpRY0b5vfOfvSsdTAYX2SzK41k1IYMFN4xwLiagnxnuSvD6LGuHKpqql/sZgB2t1lb5qyLSqFHIK3FSXopfVDkA2pmoJ9SlWHb4ivcc1msAHqkpSFyDdcP+ovSCqL5uq/pD9/mjCc1cgyVlxaLATjXd6aSVIdDjCHLONBzVBuA09owzq+HDtCZXf2YXE+vV18OOCeY8WvdrBSTR2nqTpQNGRP5931cA7v0WXtdR9mSSfkCgiFUCPlWOKYuEIKigjk6SXWAIg8s3UIprIbKLQSTzRKC3omPB0noph8OQhAyMVsh2syEUDjnq41pWEHIrE090nAeaX+luRV6/ftXZVXFAHKBciflrPkbmnlqfWBwl1MDZ3ggVLx1o/vedActza3W3xiAe6jJgvyoj608gAZq0krJ9hJ2msinwm7c4W/5W6V46MpehUl/LO94twXMgwGvZA5nsbPNfAnYFE3IfWSsFFkVI3qB/ld7U7VJXD4VlI2n1Xof4Ljq1nqXAYTiQSP7sql3veiapKbae+Z2bov+ClS6CNbGe6tjOXI4q7lzGe750CDs3yvA8XxY8bpTmJ9cags9wkqG5gqQBWlRnen7t+kPHYroaI9GqjAdRlKY+7W13RE7H2SDZGRdQBNKB08a2n/6iD9kSTN4I8ilTBfxuie+nNJ1L8xVHFUEnRwwj/PhCr3n9oPkEsNsvoHgpdLkvDPGS9ZgWZoR4CGbPYeVZ5zC9gLA6/WdAN3ONimZOwrm8ckydnNEIGVqjtmWhgeL++04hcg14JpcfBCYz5QRidR+8BycUM9oEIhVDi3bV0kdG8Ys8Hhsp85yFTsxKAPZhXXFHtd9Xwn9IbgFFofpQGwaWu1QTtI/NTpQMOtHMRNPcjL7c+qLV3ZPmVntZJKag+N2mL1MAdErbiGVRpgJ6h+JGKsNKOeO/ZGGPzHuTSitNS5YmIhRxRgCVocRt0QvC5K4qK/FQ4i//o+aI2YNdf9fqrysN77YNp+mJZ/+bzENFxnoYIdz4k151NkuMC4oMXjS84KNn3j173zLpCQuXvOi+e1aIeAeAplGAy8EIbMEOu5AP81r7nzdkGXRq9qfZE9R6AQ1+8XjPeX4TmAeRTaQp/D1liGecFL7kYWV1QWv0PulKvGHsRRRXM7l4et9H9Dz6t80ocCEkpQ0Hd0elTi5MYHTxYYjMrSLYemJEsi+PmLJOoRWXSMtxWQ6J6cEREKuesRTdsVeNAropgrucIqSw376Khq0t9CJ0/rxoZIMSkvo2jqlP7eO9IBKGs4pZyPYgQnBZj/8Ghx3utIYKMXNJ6f0Hj4io6Lk5l320Dep7z4qTIrQJNP9r++Vy1RxyUDLH4+3t1F8tv+5UjWtr3zsej13o3UG3tjdnAIjrw+UKi0N++N4Ql3K603MX1rRs+SlFcN84xqKmalVnpdgQSD9dpoz3dgareoy59j6venyXhzIXFKkoFOSo2nzfCWRSg3SCjU9Y0h2M0MtpqTSJFIR1z+m/yXlYtHLNy6h3lYIa+9CDVFi4fVUZWZHrU/ZyhZinAnC3WLfSgsi7Rm9Ew1EYLSOIQAil/U77aVQ2f9f7NMpPJT1VZRi1UslzpAwMHF5EVPUqcdsA52+pNsg/VU2GaWIWOcoWuDkNMKVhHS21hRgm49oDVlUz4nIhFQyVJapaN5Nwm9SnlRFxlXj1nVn3dYLWElYdU9BeHc64xuQAzDa3RcBSDFKwV6FT94p2ttruD22DJA0nRKoMy9/75KhnWM8t5xFK/jdMvEj39Ktc+GIMXGhn7KoyEu6GCiqrmUG8EUzyWdF0dvYgjIETbY72fnEutjdtolAce6uYOUk9HbiVFu/I4KMdPcli0WfWL9CgCpTm6L5VrV0jlA5ppUfZ79WEVGq8UjD1Z6h/RWYVv5GjYwYCIrNIzoUhaeDvHrBYLpW15lNeJ+iU2q70MzDFf2feG0BBXpx4kPKG13yx1kTpXkVM294+pfGQTyfsrzRxus+r/h3BFD+t+YczPKhvKaah9+2jkEUytPJqwOq2fW3B8T01++nvOg4/EvtxGhqO8kupKyDD43sXlZENLwFoLUAcNaEK4jQzM37nZZh0ByjGKuOWYQhqBO7buIDmc1Ry701DvyWliGawwSVF4NC+BPAIjukPk7gVQJdulyd5AHhjKuuXowBhSPuVCcN8gB8SURZGFRVJoWramWK2MvuhGwQHQjeb1O5pXclZxfO4Zog3vuRYZDxxe10eSS1GpFoL9/L2uogyOLmDzn9GRyR1ohB7kfP1qR5jGyhj/G+yRCV7zOJQGkgtoe0IRjyr7S/Gqg96zPIV0QvoIKqdTh12TzcVrOTSN3GweKVdSGHiqaFF7K76nn6yCQyldB++LpX8ndihR1vODbvjiD4Xu+DS2n9vozWudglrVIYOMuizlaBQac0tO1Uy2PT8gLmQ3HR2a/TagWoT1fBXjbqVxP+cZ6BB3QxP/bScHYZtt1zStwq21wYF7G8GZrljF4rP5zcbHhphHGoDOEanPSDLU2JqKTVDuTdX/N6+S2Clee/n9Pqr4lBFQni1HKQPvf+fxNfsVvSrKcV9/MeVCr9lrS2zKvxYwrZ2ZHK/GD/z7Ya/U46e/3iVR3w1Q5s4U4+lnAEnT4iU+SiRmhhVP7dmRnlly3ACs0qWe0YEiFA91ba3hnmWSRKQKCE1QU4TXg3ibO1MKibY32UXZu/Yo244j3jW0JyfMlc5aC+O0J7l+OhC5jSbVzUYT+zrsaM7jqnYFoANZrfV2sAhjAFpwULhF1NUXU6OCXEaVgSU9TwDTfObOoTnwZVUDUxlMouTDmj2B+oBRuZAuY5UstHgEqS6TBD7r0w2fCMUJ0dAVgmMWJvYh1Og80yFPkEVn7mo69IHsOzP2JsJyKw51SBg1iwvIrsYYX0vpRRnD3RtuPmGq48M6wkY8nFzOtATexrkJ03p/3WYtie422CNNyH2RLuQo1AUqJ4YE7FUmo67aXHXbW4ok3H9+Hd4MVGSabVhgDb4QGOv2yqc1co6fA5k1RdvlrFcTYrkeYBbBrAuMJQg6uY6uesSDMMCSsurDUfRhbOcTAKp5T2gYfalOVYvy4J2EGH7bbyG1ss8b7tnroisE6rWCFR/fZ0IFgFzbfrGd8XZ00e4kukcGXeXQ5K4OTo5ysmNH9MiFTM5+WT/1Y1TGloN4dTUjjnWlQfR+9U3uQIkK424kqWbLvs9VmhdTCXmnY3Ojh9F/u1csdB2WzK75Q1DOHO6v6oUTArAHw8nUG2DHEI7zkPahcLYbd+TSf3FA/sRQ55wVrC17UiVlz49QfiW2PHU7ulIMHtyeI9odl1llwiZ2jxIfeZP6OVA4VOgCxnSL/RGpg976BhnhNkY+dKcvYAm0StcFfbn6O+3gS2g93DTcJfnSBomKel2xFX06RNr0NgA/dQB8J7H4rhmjJDaXDoTSLjUjxfHvrArV/ABsYMy/eh0MxtS0xuq140qiIlMfxtYZFOFeqZaawvLkmyDS2Jr/MnOkF75TKlE8xKvWVYIq27MwNo8mZPqUA5G9aT90+HhdgNI5DQBKpc7Np5XTGJJyQ9PmitCvz7u1LGnJtE3zUPj1HgAsDmQ7ZqE/cDYFjtQfSt/Vd1WeCyKoq0GMiCnOggOl6UKkWZY1I8OcOWlFk2gDaGNWyTR1E1U9RIDDYSiPNrOGiX3wjOdhPcVTqSdAaEYPL3bXJ6plWamAIeKrHcNZvoWpnMv8L9WYtmrjspjqPiimr/1uTtLBiHZaW1glyH/qT5SP98Ka4dcY/qR+QroT15UJWxlosO7I3VH2YP8b2qu3RocrAH+RQD4af2SoIkTZpavcWVA08r3nk3B2gxracHw+OcyKvjVAd8xPdL9GbEIMsI0YjO3kNvsGcUHq4ByOjR6O6Lqe6kNidO2IrXmi8dTdp3kohJUWAR1tI6rCssf/VyXDx2xH0amQsW9G/EYGhXv7+gFwwG/rX2IBSaGaPp9Saa0zqxKaJBbBiVc2S6yIfRAh3ZFoAHBojc7HetOBWu9lUvRW2cBGrkHnY4XasgAAIABJREFUUMuxSXmllgo6bW9ae2xCvwqgOy2qvpIJADkLDq2GrV2+YrRV3t/zHLhJiYQlmWTm5LGefV0fF6WRhRpgfFSqI0mxoDM4z5B1ar3muD6xblUtzkidSD07Ck4hq7uzgMMuCSl6ZjyI/KHz8F+vV23cQI+CzwUbRxPXQQIWO76HwiC1hqPluTUkfdFYZYCUfMdCYPGC51WQOBaG/aGTWS1L3vyCFI9kzFGEplR3xYzyM9Ox1yFV5NHREfeQAM7GOvaHxF3OiGVns0rXIiVSUxXnmHPK9AwiHU8oTEQBWE2Y1r78mkrOJNMMIsjjcOjnAZCats5ZlWYhpJhPB5Rcxb/5KfnWerb9HNoHpkM2PhSK6rPZQI1HrBSweqfYZnA6dao8zyY9wDDmC+vZZesORNiaFjl4ntS2sUIskqKDQVSp5RE8ZJOyX9qBsx9KqXb/itCruBYi6IyHQrTRWQSQxaFk2nSvg3P2YRzJVkcXfVCByu5h+HVgAljVp6H8V5C7eiWuX1Gh+AXm9Vp8HhQJgPL54euUFx1UoCWhrR5Nv6/LXBt6OXjFwdMoqO/hYMRIEU095IfI4P460M7TlyyV8rA8sJSbyF1Cq/4Gfi0ezig4cmGgCK73v0oMx1mk1ar81VA8s/ozaiNvaPKVzboNrcqB2c4LQPfF7GoP29Fbnq4ctJBPUquCDOpEnOc8OjXrjtJGhCSqlWa2UWkOBAoRwIHkyMTx8YsXKjCrz3lvWK2g0v5NpOrqDmg5O2unv9p+hVRbhfxL8i4+iBF4ePejlAkX6ZmwHj+YvR6rUoZjCtvpyCCeohWRKJ4OfB0jX9bd3Ojfsz4/2bf9KUWHVZUnNS5BHaUh3i/7fP4mYMHhQLTJKDVq33DGWaJ7WhwL76kye6GXiLfOXCVKxekd06Kw04idc253YSRPfmkUmm0+WH5YSWDtaePJlOx6r7G0FZHRRtLvncC/5+77OfV0aJQCeBmxEEomHI4lPrBhWZCXqe5RGFmNzIKf5nSaCfW0lAMUzK+uPJUPd+ehUpESeg1j3w17UMIoEUahIKQ6E89/a2CLWHsHMA7lYK1zz+DgvSZAkV7d5UojUPm4Fnt26dit1tbEbbClWYffbSBYlkNqAppSqwvnsJzWAvSgn1MJbNwfTn+yo2+BjsdH9Z/8RkFCReVU3DU64KEtiKuxRp5uJSbsA4dyHAiml3oelvMD7NVBwkwc0MEx9brU8+8ZImUn2XyKI56bt/fVswsF1mpQKZnoveg9wa7s1S+XhkOrp9QhgT1rlH+cQ5Hqx3jXK3L/rbN0VMIyF4Z9Nq/TERdbkS2kZ/ZZ6NU8p4+ZVRqhU9Doc4gtfbrPoMo9lAkfi6mynhp7wI0UYVQbsTX6Zcf09mKQfXJBNVhle8vMxT6U6MEmkqVWjfmpKAGx4YSrIQ3/uzdHHYX1POx5GBcjMLtBzWBHLb0cWfUxlFS9VG02duNNHVSWbW1HvzJ2DgTS6EEZcufCNdfA9TXsMe6VUx+pQybgSvvefSC0uaoymflR/mOLO6yc35jdjyJhWTmAnW7qIyAWJ6vz3wA0pX1ef/VnUZ67nclEanwdUzsfA47SUDTq9BIfFfr4BPBwalR1uo45t80xJaiGKWupdl8qBY2MA6e5AV3JGtUqHs+7golWTelXkhA9q2uUnsdKiM+Rw3LfLee5bvg8qj2Z7P1QQUBVtmydkQ6tkMa4qLi1gYyfKqeuGzZYiVE6nah0C2y75+hFzQftM5hE932OSihY7esgSq2mz3bH8+QEA0mOKKlTmbmWlZafZSxJdNm4VTl3wctcJR1uIk7Rn9F2ra/WuCvd0O3N+tkuufak5d1mLuIohErUH8D3ksBIz1cde0b4tBegB7IkKDW+kKnmnmyoDRuA1zRrmCHyXCzryLmrN2TQ558WK5kdTUpWqjwuAEQgngrPEgzti5LHLJ5iaTpYRq/7eQgFJXt83L9zGQCNBL3Wmq+474dQAGBUE3HmO1r1wFrB9UaX1JQwH+4mJL0vHUQ9Gy/OJsRXiVgX82qmAsCyYv1yO9N1/91pVAvZjC3mXW7lXTXiHsapoyjUpnUUIdhEMatIHRSZriwRoceVgev+7kFKneoiO3WVnaXSZxL0+xtENma8o1fRfuthlEqU/QolYaNom0TkTInqxh8kHLrQC+2smRGIwFdVw2qU4pDCtu+zuQqzJB3n+CTq3t3OFXgWZnVNZhtfCVLu6lCTUix5wAlPf3XAIVlitf27pvbsu0uu5yg9oAgsNcDs6+PEWQTS155TkIu9Gz/He2kewWonV85bVYxongGaF4GFwVuikotTk55Z8eBzgE4OJAcdRqUqED1nYgumxB2AQ4J3JaGeYdgnbbJQUyxNZbp6ApLmXehgbI5li8gKRa3+3q/cWQ46HrbdfHazGL1AHzTBcQSQnGReWoIq0SUrLSpLa2JYM1ckzfz6q/cskoeH49w0HiDW3em5eKgSNe6DpPKmTsdWR8b+bEynVP1qnmHxmkbddxEPNS+HAvlAv7I9ACSpFxXDScS0yUgJwSKoHRm5HWYGb6Bf5RzURXqUJnuiFa9vENKVSA+qdgCHg4mN0nL9emaDdYt+cTS0KXKE6inZvSsHiV8kEdbz3UrTHaQ5iCdLTdyOwtgrZHV37KyuzImqATujDTpC+bg4Wu3qxR2DEdDt2EzAlN8bVYHXfzBysW9ANXxGbndNKrr4+nlwDWDHnQPgjdZWA1ZbzuoVNdTbEnz2grx1K3vPUkBNtDKMfu4ujUqXMD5R8GunTzKsnnlhhURKE0HSzI3l0skIIvFTcRvlKUgG2gV4sJ9jMiX4QZ2zF4roz1ICHrV9kYllJHVdYdrqAy3UVLMdeMWhz+ZAarhPSZO3uEkORBB+z5gAtQ4Gr5wce9hswVcpSAfUpQjCVXe1cyfG/Ox/cwH5TDvxPjsnVTHrtVXVxVBr4UoHKuXwBHmHfZ2iJrPvzl8isqzXbfulbdW/lftbk4vj9YfPVCK7ruRxnUqMZ6gZH/UsWqPiw157/5DVT9IKzz6uAPasGO1xTXYr7c05Z6M/o5yTnjeDfTvbVrSeyN9cRN3INyuItopX9gu0JD3BMnsh0LnWbfb+4kNIdILOKTu6Pz89hFflql0OwkYgDqRx1gF2Sa2mATG/588KltasTr627sgQkuF7/IbkfAb6xxTBp/JmBDJ1NcGeiGRks7fXLdgNzR04tAK620Mk1E5FHBGB5ICgvoioB4t4d7f2XSwSHHHR2YbLHhDC5BQbTWfnQl8v7FkdlY7t29bPMnbuCLbuDiqFrlhqzYosTQ2ztAox+aoepCKWDK4ioDp+gRq6LIk5YD07JFHVl7i/63fXzQnq5Xw1J2HPh6i1XfkFHM7716QposWucJG4DXxV+vB8semKv09+Ya3t6EMTwxjw6rCzbAxwwI40NTXsOJ/NCalCEziGVz8/rXLsy4qXWgaCwYx8CnutdDm49q+rfvD+XEh2rqrjs3kPr25sBUu+hhBrpyBMI2BqNGOq5gocC6VtdGT80Fm/oBEIvSaEn04HNYd5GifyaLFghkDpBbpKYgbLSfhPtaQ2/aiaOAfcGF6dr5qNmgHR7eU1lLXbzU1qw/qwcUDOPXyH3s4OVCBew1S9IDFomh3KmQzjhfUIrcxeDNgoLp1scdBJVTSoyKk24jOF8lFj702qOjY+aZKVpLWbP9gbC+bCkYv8ColXb0aOjLcatQo+Kv3STIKk4s7Kq9T7j4oWFd01m+BpLYa583dmpzGa0QDzKvHyEIccala/R+LVB97HJ6C90cGwEpX5+ESsn301w9j6mcwq/fW80pReRKP1rt5zEK7//6Vn8HKYzisQMD661V7VmBbV0X79VylVM0N+2285pJr1OjSFS81jqa7SUcOC6AAGkYDrWgsjgtVs17HXV+skjoZeGcM0g+LZ/IYPIGvKmPuFtSqNb97NKoBW2mSAV3Of0A/IN+2uYdMS/kLJp/2qMVOBznbiCQCYyvtFQkHEHCrq2pCkVo1Um4CREKpJrNR4+i30KEUeczBJY5uQOXoPCJMTnErEHE+vv1lebBTQG2Bsp75huo/TKtc2PSOjTLRAphjfCI3LR+XdQEdJtIMoDsO40cELZhJri1igPhi19AtuGzQxytn4pNRtqwfVo6ADTqfJfH/fXFa8xbC50QUu3sjmAA5DTTVD8ZKdCgXlDJmnSk2q3Hr1/AkdKg5CkdHRSBM/5FqsUWYJgFDkpLQZB5/jfYDHPrRUvv4Xo/z53BJt7RLsaNJyox60fUKEHp1upXGF5371PWjkHG20TIp8E4nwnqaVi7n9U7S+qcUf0NxNVZv0nHUGWHIdsSN3k6s1z+JEQU5H7Uw3PMH9If+2Kg0MtZLbQAYnZOnkRs0/EaeocvLOBBLQuEiOc9jVO+z2BxAcNDpOZKyc/YV4kEqjTGVUen8e8FRDWUtpWe9n1IsMjuIyuAU9neYYKmJvOTG08XJM4kwk7OlDvRvOFKHqdQ9Jql4pC06LU0g2S0lA5RADngXV6AxqtVlEaq8vjbyco642eFANPhW9tKk2xD6jc8xE8QRAYt3/Ogxbnp9OmMgpl/pqrkYiMjB9tpI017OqdV+HUNAWNGykiL/NcCtU7/SI6ZYitw6FeXM2YK6r55eKszUriq78vX2SObUbqPkRuhibKZd4EqE2aSDqm/j1ua3nv652OFK8bkk+10L2FqtneIJ7tTubq0riJhQTOOeSqudCvRGbf9jPrv3ZjX7ZP+eH7YsD2BWvminSIxcgcld8F3awpU4m14NdbTxmlIjEZwqrc7Zb4aUAfZCNKudWcKrKZMeEMgBL09vGBaunMMJpEmVdbViVAxOi01yKeMuqWPj85GivbPienDNR5Tm9LhtksEtmloLTN6HnR6+RdRPVNmizC7DtNWuRjluzIiHiTxDM/aOdD7KgKIwlYUcZgYYCZ8Li6fJdG7wV8VO/o7r7uz6LUh8f/PxyrmUULiEXN2zMfyCp7VB0VGlVh9+HE+JS24JRbf65oKvndK9JcN3qar/6WfjnEX31lxUS0sEPpnmQc5ztIItUHgV7nQcuDWN8Msdlrwf3ttAh9oAfn4giriAtSzU5kVvBVm3Ws2zF4XZeNHrai1Klup/23euytTvbttSsWOpHHnaog5mtC5JDO9XAIt2PVFONXnsA0Ow9V2Oi8S5WKF0BADuGCmmPucYlsVZpHB0cnUHa7YL7BwJq6PysPceoz2IkYptbWcicbfOBN9TL0qMGnBeQZwJeF1mH1ostAn27nomINvRVlwysQI3VKx8Xx+1WksDaQ4Mb9IA7ymQuXspDQdJ81WWvFk0WZWj0XUGkyv8rt1VLN1h+rUhxXF7sFCrlhchbGpuCz6Fx8EybBG/jgSYP9TWKnExdcw9W5ZjY4+uQURJrLopI2Z5dkQu6BhFIiB/t/FNa/ATgWza8vbZEX3kQSAkNx+vIQigKte+vN4VaBUOhPVKpiyRdcDS9Pm+lenLK0UaaUQa/UxzeRRt1eANP76+a2jJLDuwWyHxYLUq+x+qLjJQqAgks9ZfM3eJuUe5ycKRcE7RAqS3r2kUkm8l4FWaXR0GIDaDLlkINtLM0NjnGEaHXTftVN6U0NKpyUQ9ijj0HJfhaLFk+urZg8czssqb9W4NfsOlLexzI5ouUhtWz0S7rf4jM6rOt/Ko167mvlB4E0zppH/DsZ4mtdykno8CQ/fn0R+p0CAHLfrunBLQLIpKgPihDFOwmkdQeXJ6vWmpdUlq/ID6/Fngwcv9+I1Aeq50+R9D3ZT3YkmDjw5tKhSzfqE7u8niM+CKa+nVByGdVjj0vftU9FiIk5Tmd3lgb64q0x0Ham1lOqVSNYqPrc26tg4yx3mvXyJXz0eCk+EymOTj0Bazn78hFMkxEYO9N7u+b9ygBbhrMRg1c5V6pBApGULMS6Cg9AEmvLpORuTdz6nn20GNAZWVjNN+/D7622fFvivtch7uNdGz0dHym+j3ba25CBRvai4TX2op87ueD0lk/UBN2S3qvJe1Xdqs9PGxSa1p/H0pkiPSWQ5PcfxxrvMc+dKu8bLSrL9X4KNJxsOy9CW3HYeWNpPsSrl4DldA5b1bE/+F06zNtrgbNTeHXawEoZKYmTZ7naXCSnmJDiRRMhNpgE0xttuZFOIqF91Z5HRAQ5T1dmgtzBBzDrmaStWXK5yXLrjFvpVCTsZ8GBlDmrKpH+Trmne+WKRudjPOZCrZuyXePdQ8wNRlkpdH3YNS/NZtAzL23gZt5DW3pA0/tCMuRhc7q8ynPl6y+yqNEbLU70E1jmeQH1ul0VcIaRAvMgfN0mLy41zSNPaoaARDCP+04VAoehOKg4nH4tfkjQVKolBythUkYhyJv+OqtPAx+b4t7xIUZvJ95ax34X64agNOp5UJXi2h/oPPrDtHkWAUqcaXJcNMVBXQYPNLbrst2aro17ZepJmhz3ge/Zk24TSpOt3Mr+y376jGK/W6551z2zeix39+caQnYp2KVImrV234VuNHrVbf5PUg8bZPwCzUeLxUmepgOsAsLmrqeuae29efV+AI5DfrKNMtphpRSU+Uk5Kpypl2H0dTyZOx2cX34Pky6iAWSaQwa6mDb62rvDjmi9mgojKSoc4iCYEw/6dB0KQxjOGpWwjfk9IqwpAIuDJpNmblYdou6CAb/H1tvHvXrVZUJPvu87++7Q+6QOSEJIQkZmMKYIDLIrKg4IrjQ6kIEbUtbW5fDcqiybLvXqraqLBtX21bp6lXLLqu0RaVRVBQVcACDIBABgQwkhCQQMid3+L7vfc/uP/bz7H1+d9VlheTe+/ve33nP2WcPz3723qLtRsOUyCTEd+u/I0MjtNvZ6n4f02aDdV2ZqSCwlXUoe7C2g3Wp9mjh9i3ITkneYZsNuhd3pGMPfT0dF9v3mC0JMhzahEsuPQfH5wW33HWK3K0qcmqtAVh4PhG3nnXsKK69/Bg+d/v9ePT0giaQt7G2wqowSmEV3LE5eBDXXHk2Hr7vMdx9/2OI8Y8bXHvNRTj10GO468vBoYFZNDtiBmyewzjsjmg8FUZk1RAzXm3CzoGD6Os+lqUAWSRZiCxYkosO7BzCur+H1VWe75TPKMyLJi4zlXXI1zQZ1r5JWZXyjszDBpvZsK7AumqcgwxSrCVrdXRbmC2ZSNVP7CwBYaD3NUrSsT+8u4yRpfdTtVdEjYyT20BjLfBVIK68YIKdYBcuR9QOQQTCZRfTzNC6ryn3EdoH1pTd4Wxga6vzPCxbESQ2V2Cvzd5Xq5RoQ19O5SXWi8SlHFBfiwVX63AdSAcsqkq7rzBW+rW2wxme1Ug3nyfL0VhQte4SNOW0JVpEzR8NhJ7NapmyEvqdc0Ut0prrchqYD+UAXPceLDsDuoveu0uLbMQEllRAx88+guuuOAe3ffYe3P9oNNHpyy5ueOlz8GOvfzJ+5Kd+H/c8GmXxbW646upL8cqXPwOvftHl+C+//Pt459+fxllHz8LTr70YX/z8fbjry4+n4F79zGvwr3/wRfh3//q3cfM9kb669NIL8KIXXIHb/+FT+PtbH431+IpDx47jzW95Jb7hRU/EsYP7eMubfwOfvv8U3FccP/c8PO95T8ZrXvkUXHv4cbzuB38X3YAXvPy5+JE3PQ8XnnMYf/Jb78Ev/NePY0xXS0mL3SpF/qSnXI6f/J9ehmsuOYI7P/4pvPVn34Xzn3gRfvyHXoVnX3UcD975ebzlx/8Qj677OOf8Y3jOs6/A8599Ka5/ysU49+gO0B2fvOnj+Mm3fSh4K9zLc847jBuedyVufOZleMZ1F+HsI1H8dNNf/j1+/tc+gi6vxPZwwUXn4MYbrsKNz7oUT7v6fBw7HI1k//rdH8Iv/D//CDfDuu7hvIvOxdWXnY9Pf/JOPHSSmJsBL3zV8/FDr30Cvv8n/xAPnd5Hm2Zcdvl5eP7znoTnXn8JnnLleTi007C/u4vf+LV34+1/fW8ZGXoxkkGFRQkmL7uJH6zqEwGPebsAluVkAckueV2yATOMhWEie6mgTvJLT9uXXazrqVRIvQdJy5ze/Ro4kveVMhvPWvdPQFmvURHkWrxYyYDSssReBi9ExZfdVzR6+bPZzJyVMhCVs05Xhr9TcktW3cC0IrGDzmIbuZuAQgfkc/K7mDFIF90qhRbuULR2j+49CxVKeBQT0VtYeDuhLIIUpbRsaxt4i59rqnHwmtjUbIpwA0CV21sqyue//Ln4ibfciEvOO4T/+st/gP/r3XegTRNe9rXPx898zw144NZbcWLZ4CUveyqufeK5+IrnX4HLLjiEf/rUfbjwwsPYP214+o3X46f+xQtx5ROO4O/e+QH8xK//A3rfx/O+6jn4uR96CQ7vPoj7Hpvx8lddj2/8mmvwlCvOxTnHD+AX7/ocPnzbCUzzQTzjWVfju9/0Apy9+xDe/7H78JWXLFjOOhdf89wn4NnPugQveNalWE+ewAN7M3aWE2g7B/Etb3wl3vyay/HOP/00vvVbrsctdz6Cpz7lMtxx+304vZAW7UqlRrg1TYfwrK98Gv7199+ID7zv0zh01tPw2Vvuw3Ne+jz8+FtfhM/8/T/h1mNPw8O33IsrnvlkfP2rno4XPucJ2H3kUfztTbfhP/7HT+KLD5zEq7/1xXj1FefExKsDM65/7pPxda+4Dl9x/UV47IGH8IGbbsev/MXN+NKDJ/HaN74Cz33SuZjajHkz4dnPvwZf94qn4oanno9Hvvwg/uamO/CeP/kYHnh0H2948ytx1RPPRjPDfOgQXvGq5+N7vv3ZuOicHfz6L7wd//n9X0SbZ3zNN30lfvxNz8Y9n/gn7OEAvu7rn45Xv+xaXPfEI7jztnvxgQ99Fm//f+/HiWXGj/3E1+KJF54Fs4azjh7CpRfs4PbPPYTFAeEnTelEl2vPvxsZpThDflt1AY9QQ/JLRTDJWjMTwV9Nd45ZEmOFdWT2ALc1w4+Q44lhCKkLAGpotiURLSMBhXPKJEb8ntmmpMefgRe1NmOB+ey+BFREcoY4Dk7euDRbhBmWl1SXL7IQw3wQOkierugMgUmafJ0OmDWi9BXnQWQcMMvhAooKghVYpMpVAWA+rE2fHcOoWFfPTUpoUS54MjiBiy84iD/+45vxhtc9Ex+4+R5sDh7Am976CrzhJZcBs+FvPvh5fPcPfj1e/4rL8amP3Ip3v/OD+JuP3IOzrrkOv/ncC/CcV38FfuilV+Ij7/skjhx7Gv76I6Fsvvk7Xorv++ZrYBvDB99zC776jS/Dd33NpXjHO27C77z7IH7hf7wO7//Y/Th8/Bje/F1fhde/+kp86M9uws+/6x786i99K3YfehT/6ZffgHnvFP7sLz6Bf/NvPoKbb3kEP/bzr8chm/Dvf/Gf4VmXH8TP/uwf4cWvfxUOG/Cd3/daHLNT+MEf/k189gGBWEyZQpwXx4tvvBy/8St/DL/qenzLxQew89Ln4psuO4a3/5f34aYHj+A/vPYw7rBn4Fe//hg+9oFP4ud/7ndx860PYZ/9OY9efDFe8fwn4B/+/EP4zje9BC99wZW4+tKz8Fd/8XH8q3/1V/jHWx/CQgLW8UsvxStuuBDv//9uw3e95WV46QuuwlUXH8Sfv/vj+Ol/+V584vaHowq0bXDelU/EV11/HO/67RN46/e+HC95/hW45KjhD/7yM/jql12Fmz71JWwOHcD3ft+r8Y1fcTFsMrz/A3fi+3/ka/Ha55yL//b2D+P/+He34I4vPkaxmHDjq27AlUdXvHfvEH7iR78WL7zhcvT778O/+PHfw5dOsXwcQXOOMDiwhqhNQl2mtN4VZiT5i+Fla0oJKy07gOdmULW1j39vxX1Jz0DhhIy18ezk3fQ1MnLucN/P+5vhKnumyiCHt7KwyhsF8pIJ3dl7hsrD5r6usLWmqOtXgU9cbCK/hezHC2pgzpxKoytl5wuHuEwR3mwmov0dQIf1dSjUGnAI9uDMyVZMm8V8UgKL2gCuNbntBBc79qPG3xZEF2vOi2RNhzpsC+fYYg+2hnf+1vvxph9+He7+2Kdx4Ior8ev/64vR7r8HP/zTf4x//7bX4Q3//GW4+cOfwXd+x6/gjgfCLbU2480vfjKwOYSLzlrwv/zUb+PoM56Jp997N75kx/Bv/+1rcNWhU/jpn3kHfuBnvgWv+KavxBWf/jx+9Ef/Gz525yl821tfi1s/fS++4mtuxHd/+3Nx32dvw/e+5T/h03c/hiPnXoC/u+kW3P2Zu/Dnf307PnfvoyH3bcbRiy/Cjdeei4MnJ3zwnTfhf/ujT+HB0w0XPP1ObL7c8d6/+ixuuvke7C09LSKA6Ko1hQe3rnv45V98BwDHje08/OV79/C3f/NZvPfvbsOJPcPVz7oO7/vrz+CmD34G77/pC7j/0ZNbcmHWcOll5+G8wzOe94Kn4MAn78Zv/Nof4QMf/QJO7tcF8R4Typ70pPNwfKfhK1/yFNx88x349f/znfjgx+7GqX15fyVn11xzEQ5Nhhe/9Fp8/ON34Fff9g588GP34C0/8Z247cP/hGPXXoP/+60vwd5dd+BH/uW78B/e9ga86XtejQ9/4Ga88bt/H3c9tFuGjjL29Osuxs6Bg3jNq67Bhz98G372p9+Pm2/5MlYOulbxnRicfd3DNB3A6qcr89eX6IC2emFxZBcrjd9aMDODgd2rbQAWqBtVFL1VZq7aW0aa2QGIEiAl0rGbBnYsTOtkSdc9rh6zY0MgfbciACiFK1BarQtDUOLVnnHj9zxom8vO6e7ZdafSfpaTmROnII4QreEH9t2QRkoGGbWktQ2xgR29QimbrF/YSQ+hs5QXXs/IilWy2Vb1teQ65/kwluVE/pyIRY3dpMM1Y6dwZja0lrAGawqSNukn//d/jq996lHc/+VH8Afv+Hv83ns+g5PLhMsuPwc764K7vvhvOtWkAAAgAElEQVQ49vaXQbECT3/edTh04kHcfNuj2Fv28c/+52/C977qiXjwgUfxV3/xCfzn3/0HPHTKceETjuPsHcdd957Gyd1TMDT80M+9Ea977nn4/B1fxO/8zofw7g/cjj1mtpIHkLUxLfd2PriDV77oKnz4ps/iSw8+Et2ysjBIghc4UbIVKfCTSHY8t5UYTu+7EAdEZc/VA0EzL1ipqgzMNOH40QPYPXkCp/aGlotUKpVCbIB1nHP8CHZP7+Hk6Rqnl+48f0UqHDh+ZINTp07j9C7bAXjDz73tu/HSKw7g/vsexjt//8N4x1/ehlNLw+VXnAecegxf+NJjWH3isU4AwmA0mzHvNBw5tIPHHz+Jvf11+F5mrZKTAdTQaGDk4Ej+wlXfGbzv8myTh0QlkWDl1sBqYJoPYdk/wfOI/VyWk9HvBC0n1U2aL2tN8CiU+hXuNN5frROQUT2AvpyKmampnETG1GeZNJAht4b19G0P2zNueMsDmC89t8qS4zVzkKt7doTa+nVGDjprAMaWbszlmzWsy27MeZQld0/gCLlYgqzrLkR/zs5Ek5RJpbaA6jAldt94KOv+KajvoADOiU1Mi8oseiyBH6UG+4Jj556N84813H/f43j0VHxWjD6tR30vQiBU7kx6uK84dOQwLr3wCB68/2E89BhnlAz8iqJfG46fexRnH1rxxS+dwN5aCi4+p9EGVSg1CmF2Per7UMu7LIIji6+r8hDq6WAVOwukpsD0vubnJjJ1xR7UBRqH/Va/iIa+no5O4KM3kVTxUSFw46RszSDgWudx5vO1v33dw7kXXoTzj21wz9334uRelQaEEzGka9ljI3klBNZjXORaYbF7rlM/qxGF4eKzFZ9GdjryEmuPIUNGZdFYmFZd5LS+Ch1C6W4ovyVDy/6JGEok5ipUMj4C/cLZNPuUmZHh7tQ9FSP1dCgL1rboDqspk3CNQgYmLKdueXh2d1O6ZqzMswQLO2lfoulWNyJtfEzcnlKBqMw3PhteRlywUiTqCm4wpsyiuEdt5Hn9UF2ipLwUW40cgJWKiAVv3gPY1tuydBuuwwlrE0K3CzalpEVoiVA/+uDDeOQBVnMS74gCNQ3vNb4bwy/FrKj479RjJ3DrYyegX53uqSmebJaY0CMPPIKH8xl7WWAFGNAs2YkSFni5oK7L7Z09UtlblLsUOJAFg1JnK8Um5dbLi6gLrqx/kfG0zwL8RtnQRdA/oQTkfTDsM7Vl5L4rRemRkUiF0lc09p5QkV/c42DwPvLgI3jkAcey7AUdPS29zp5hRxYBNgSvMhRDNuyR0oRo35LfSrf2dY9NYHQGDWD7w8A1iO3BWZe0pEHKjIhCkD5afRpFYQvE1NIwer50yJQGIjlCiVB+xYK2Zinj5QHVyMQ0cIn3dZZ18F8WTO2RCBctDhxR4xpBGVbfz8G3ysWGB6nUjuisJAQZ32WtA+7QQB/BQGt6CX3ZHX6ob2tMNmUxVMdhAUXqVZi8C9SlUep02T/BuCueHZyQPbgdRBS88XkT52iiKNPJM0hBbEUA4kULYTeI712jFlGl5Kmcelk3eQJ5WRgKKBvhBV5p3yPUAqLHQbxPlCBEvUNq/i2MKXAZ9eBMUMvXHI/nOQ+G/TN8TXDLLEblrftK1+1xIlZHX6VYqkgpq2SpWFcwJYuWz9cMjqx+VOGe91SQou1vGRvNbKUS7Jo839SyLpQ0GjN3Ls92P0hFzn4m1hBtHRjPsx6l+oRO6UGlNzpU/4LgnvOSrezhEf0n9gdj07KUPWgDu1RGahMZircLpJQS43PhUa2rYrSohGZHb9ICYuEL4MGydazpHfKloHsceyyPgqlXZ6Ffp9xLHmDZsEdeHJgNUshpCGU3o00m92xiF5/irseiEr8gJdr459LfJRDxE3KT5VomDVYdoXtof7OBHSkCC7Vma3O21g9S1zgYV9YDKEq6cZMNYJGRsibN5iQDVc0HqeMkgOl9RC3P6VJ8v2pDb7nuVFi0QPGsKTW9CuJCUELpJlg0ZoAgWq9xehVj51oBxtL+5AEwrRUHPdMIDeFhZxGcRT2MhiCr/R16pYrLTS2vTmX/47RxKeeiUA+dy8xy3yN1LZ5F7WXMC1HzmU3+WVj0+phi+XCqxMJl6s+ALFSTcjcgmtgyk0F3PKZZFv4GIEpPulr5od5HTIHEg0imgifNPBrsrvyZYRLbaCzkh1k9v2UBmLwsiy1j57Y4U+5hI5mMDZhi/9XyUB6C9nXE3MLbyCI9enywgDJzP9kjI4x/RQvQ/eIE7IAQIrxqNqEhL2oBS1HNuW3xkO69rJJAT6VWGMLkz3hakVCi/FnNXWC4U+kaeQXjRTLGXR2aEq2KzUYmmyykvAqnK+c9BqbIjSz1XBWBSvv2Xsqxr7uoeHLJdStlFd4BLY7XhDbTYUjIE5FuQwilPDfombXcZ+1dzGQ902JQQWs/UxRQHsn4jq46C15Mdgsr1xyoWZuhBMwVFk65/irUGwQPShHWDA0fZCKWHK6uzmUkKamXZBtkrPaKsbPOiHTr7feyrFT1tKJetHcXz0EWUhog9rhrVi586yy0bgA1s6R3VD+Hnvuf/TGFKem85RmRGwGgvC/ekWJFKvSSfNLo5N1gdbL29cywz0p+fV3Tu60eJZ5nI08ilS1qWl4qCq476Ao2yBBSibD5TQeMHANqor6OCHVZaep8wHtx/+FpmeGOFaHZOhWGrKWzhT28M4ZDKgsA0aRHz/OI7Ve5rETxAwDdh4EsUBjQF/QmFxfJ+AzBWslaY+m58uTuqXjMkc1apEnVIyG6Jh0ogeCaKQohnwn0SfC2lWw2pTU1b9FIA6M1HqxOXo41LYGsdvBAmGnKwj2nFZyom1fA2LSVl1wuJ1aGArw4cZuCgRsNf4TXAN7345M9en5GmBqjKbtCRJb8u3dOfmARHtmP6heRACNVTpxtlyTFFRjmV6xgpk0Vj6LUE6GPVvgtKjOlEJlhAQxY9wN45KVSxbQUaAfDK4+LlXwCXvwVZGbybk7KAskDdQQ4mG67x+xZFGAsb3ldQ04z2yawX1SDFq32uqJr4jOt1TAshRxBMNxJ2XHj6ETvqUBVOOmkewvw1jpBJdLmHXo2MiADhpinYqnk4I5ZqK2IIXKT5PplOhWgJttPzRhIassGtQKJ9GXBUAtyytRU0BSLmKYdCNXO1nt0rxpz4j37Lowp3BZzDAS2OhHsFvx6lXk3XrwmrIN4BNzzWW24xFWj4jB4doVqxjb+iqlZPCePJtvBCcBV/trKmslwqi8oMFRp5jE5C6dGz2rw1Ih1gCjfJEUOCyvWoz4kivdifxqbskqRxPexNV4bs0sB6gXmNLL8ZhZoGbpF0V9mAhSjs/0b8rIEB8BgmIbBw+mly/gAyKlpg7sOy1uDznNTiBZhY0MMV5u0Ffw3FT2ozJORS2UhRaXWAKaiR4d5sY01pFheV3awYn+HZo2KkRm4dZeZEHm6CEUHTSGbeJ+4BmtQzQu/NsOO3kN+jVeomWFSE2jIk+pR7AfBAcwg9iXvja56nFsDPErkwdC2sXoVrFMqXLCoDSFDIjEilEXU5auIqG81l5H1aBzc4p2j7QnOSckoRu3kyuvAYBZFW22O/L07JlR7MacGrxgwBHVdToUyohvV0y03Wg9PSxjrpdX0lWQVUIPuo6/V8Sl6MuwgU2HM/nQPFt5Ybk7zSlr6BpkXzyFIVX2a4JDcc2ZVOqeQyUTFwYo40zPlm0oXCm8WaNL4KOClHHk+vuZ/1yBmuv3WK09OxV0XV+e38hJN7I0gi7/mcCN5X+t6OtcXhoCNaB1QOCiFoeI2lUpv4zNAa8RghIc5V9kMKtvvPfp5oBXQGQAqsvLZRhffwgvShXRadDW8Cfld+LmOwEm0FwpJhM+tKb8a+xC8EoHfQeUOYlWHLyvaxPvA+iHJk9sypKkVqveKigfPJNYfBjeK/BZ0i6RCUgyY3tRMlwCpmU7uC9pUfCdlwAqrG4BlKRUbQg6doUcZQNVaAUDzueJd58h3krLAkMSR8U80blUqs9KfOdVKWQXV2kt+HFBPA/XtDG05IdWoMBEzqG2+eBu+Dt2FsrxaoJcuqYa2FLJb1asTmjlzJAOvYABQI4Yf3DETU65G5TlCq69+Kr7ZpnAzefFBJVnWCcguYukpiCWHuiQAOqsHM61mPV1C+R/Z7yEzQnx32gujGy1PzTQAj2uRZc9zUWk4EHGqMBRd7IHNaPysQWekegOuw5DWLkNbZ0m4QFXuT18XZKs/KoecppaeRLELszIWIgau6XpLXgOsHZQVBDCDXuo4YiDORVkSSOERVyr51dmpaqMljiHPJQXci2jIzQhpNfJj+IxRaYYIEMxmk6bw1HmemSCY0WwM2mz7kmM4V9f1EiaCDPegERc5QlRcDd4b/oBaG+juyyDMzSa36WC6ofpwuaoEp6awdOFqdzjTnmYbajOCW40u+DzO24xwRn0kNMkKCLc+mquMfTHaIKBGCzzWeGh/ymrFv8UNkYtp3MQpL0TWlfAZeYANwFpxqmK+PAxZHyqX8iSGtnw2pXDp70CF17PPBGNreSVxUil0QRTSIB3PC5Bcfc23yJ93pMKhoinFGs9NcBYcGpXkLlqndDVrT0SrF8gYMTTgusTNtt7RFSZxf4L3QH5HG7IkZtkzIi7Y0KAmsy2hFJLx2w6UggfgLS5msB0d07RmtbG8D7gnoUpyCbPo3+FqWtRhtoM2VSOkmDvSgEkENCsPhfLbMuVLhcUeI8aBTRUuAoBCw5bPk7HMd0pKwFRypPNjOMzgdfA2a20tQ9JK9xrpBtmMl0YkxE39WjzvV7E4w3NNbxkM8x2Y13XPmqkjdEmMu6ixQ2rNq38CRSpdPglMvBPje/4+uloHKUUTuHRJBAiFkloJFNFl5GaJDFUxqiHjuLz2tBAmrcssAlv/h4DXRZ6muMBZ9OMeTM++5IWuS7ZBNjXxSol236Ongnpf1wFuaJnpKSVuQYxE2A7DoYbotdhJyTab0BECzQ3B6OKLAiwUXP0/UqEydtaFD3e6sKV45MqLrD0nD0EDgoeQMv4tz0HhA6nRQxgWyjLOL/fSHekCW4OtBFnpiXTnLFoaBWUMej+dF0lzSEVldu/oCGA2O6andRejUSl0hcTRDyI8Z5U3tJoKRg8BrcYUSEaT6blSNpuIfQSF28ClQXhWsSfMmKWhq9IAVUvLm5WxcHrr8Zk5wVWFTvW5yrIAllWjzabcp/jsJvbdLAczmweIn708iMfFPgj/EdIT65tb23jku5VnphXrC11VuS6d3seM7qrLiLRiaqABSAotr/0uLT1lO/z487Xv5oInNovN4bE9lt6U7x4vAz0S+kooroS0MeeS8kAVzyfANnopxBicPRuN1rYyHJU2s2lmLDeltQexlqSoC28JLUIAuMhsEso4FDV0Md5PvVfF7zoXdBA/aikoRRePtGfuFd1M7VcqDV+iWbIUliyqqUHPVOX71uAeaU5HNWHRcGqw27b4CEmZpvfTrNih8OJVaJKWeJzg61FT8Xs9vFZ5B8oadX1+Yop0cMdzIl5wFor/wzicGTJVlMaZFicj3l/PMiRQqvDa5qwBCU8DBHxDFlrKb+AD8T5rgdkmklcxRRuMpDN1TEN+f4YS1tJ4qot6KNmREgDO0z0AdexSqKHMTGa6XFwq3TXLfcvaHREWocFcU/irmWZzMMfKh4GdrtJqhvVRSie1b6dF7YrvyalIz2DB1HhQ/K7I0e9nNBjWqLO+QcxG5ellTQ0lYhQSB9QGvXLwFFhaxHT/M5amB+YOxWXqramYO8ljXZsmjVw8AFefAu1Zjy7bSmM1WvauoTS6xnoXgpm5lwpVFA1x3xtavnfsYcXNTnIW5BU6EqhNXCTPjvRkKSKuo7FUvbUNacfDPhA5d3phebm5F7WXfbBaOpc4D80j1dk3xeXCwvScVHNlzUKcOKXOe8qEMkTyPFMpQvIrzkjXJpAvs+ZnDD7sBRXH8Fx5UyG/B0q2HYC80pTgeL+uFDwVRd2vstLihIx8DvoGEH7YuHZz8Hwa16c19Noj7yX3W/dpSRna2lliImpPqfMTm1rb1UwduvZhBmsmgdAnhDFkrD4cpHEZitWVgqFgik0oa1UbhOFFQG1ukU7iSMStv8uL4tyoabhEvrVJKp7RZhvEaNvPDYrvltWri9J0ASW0aKmkfF3yXYtCixI+vl8IB8vus/U3IOo1unpv1Ig5Kd1QdiJ6eVoH7wvHDBJkXfeBvjIV2gH0PGBgSIX1pfZPSpEHmCLUS9BausxLvo+LgMbLpEvT2kwl4GgJVi+8UAK9hw5MqMvXmGmIHiVr/lydufa0lKSUqtoemk1bSjOV1ig7UhpednVLqdEVlxIspdG21lkhJbJPZ4ay7rAELFsZjLwr489HCBDgvlY0Kro4s/herSv+J2wt1j8qgqIMtOGiwysFWnvMQL3zjtFAOqR0w2BnLRDf14a7VYZmQU1BoScQsxypUVmuPHIQ6t8tXRmALemU/hsutHml35LhSddUgFziIPQAet+P1vYu9p8jJ60DVFqoC9Y1hT04DvBIofW+BtLQou4kYs1NumnxCGIEjeXZNkF4CKR4klBVFyMU1Br9LIXVwDOtlmEaXW7keun2pzIWFkTFaAJ6W7mECEFf2d8j3HnRhYMQ53kmDJk4z8IRQ4s7FXS4xxH29b6iMewCla1S4oEfRSsC9w00uU0YgKxll8KQG5MCyMxOk8WUTCgkW5L0F8JATo0z7NLPEN5XCjN+lgrdlOoWMYsXkF7h6r1KxyGDABQGg3DxXUzWyg6lwoNqlZBhrrqaJ1jua6yb6qmKwEp+M3Qbf5lKBVamkxeY77CGhVQANtxBpkiF9/Rco7qdresu5nnDv5dsyXj1fNdwBSb0DMdDXsYCTZkZ7a/B0BTPQJcwPQacsYmWmjU3BEM8SAHL/n6uQq2V1nGPbo8lzyBBMgiPGOnfLILy7YYecq9iwpbnhUo3WZuvvHkftGdq0wEoI49D5eCdPIre1aSHIBzH06nNmopzolehLJozvlyTMZpFcflesd+dJcU+KkygPCL3WqOHe5tIeJ6Z1zP5s2mVoe/W2kTLRrWK31qHmJFai23t1eh55AVN9xZUKo7sqgak4lN2JwvCqAjLiyEV2zVpTOCyPBTwvcaOU8WM1fdl6/2tdKIUsyy2a/UDJlXeX77f+O5wqKuUIQoqU2Eij2HwKhDvQBlXaF37tqaBkHwl41Ver4lDQvn1FVCWLOV3SflNhZh7yGfxlxSeOBcynr3vpvcQ/1d3yfnduo8z3C2ELzgFAW6FUmhtDsIU89GiuoKujSc/vVDg2OchVst0Ylz1JJRoKhc/V1kN8hB8RmQWFO+pv4FQaFkYfasAPZF3QhjbfIB/a8PPNoJ8jeXaYmRSwNpQSeqAYcLcZnor++GWgimyJjKMOkmH1yFhnNjVGswGCWmuUYJ0Lk0t+AVudpgHVdoE2BqiXL7LOjYCvZzMpglbXZd1SqGHsAeInRdZnNbmBCrRx/CRF6qZ7iZc1sfAojhPpSZvLGspeEmUrkuFJuuf7nD8qYrcQADOyJxVpWmwSXkRRyyA7QfCGpPXIEaowgTtw+Dh9b4HqO19Z4Mghhhx70hHpzcSCwPJfZ0DjKwUIwYrTe8m1yiPsseYShmVsvrF63FiMJLf6IqugGpicaDCMcMaQzYSuA6CI0MqhimGCZg0AnF/kNMJk3hJKl4DgCw/mACG+CvMZ7PmBtbkY4PU5katrPQbDDVjcxoQ3gku+qqLJah8+DA3hOBJ5KltOPTIdWdJLb+/2Qw39gKweOHM/ypdp8+bDZTdBktUnBvURZuGpJ4u4JjakzvechUQQ7QBvTPvP7ynNHiVavP5MLRkfYYlzUYkrjoaS0URYOz4/mFvgii0wZGrr8HZT7kOZ116ITaHD2F54G587u3vwv7poJlhmnHkistw6s7bsOzHz0+HjmLecew+En0n23wQF7/qpXjgfe/B/i4wHT0bx556Lc6+9mocOOcomjke/Nv34p4PfzqU4zkX4fJv+DocnB/H7b/1Luztzzh67XU4+ynX4PATLsR8cAd7X7wNt//uu7Hscd/bDg5feRXOfdbTYI99AZ9/z4cwHTqCNq3YeyzmvLaDx/GEl78QX/6L92BvT5kfoFJ1DjVQ1j/R04Lp4WaVJbMJ3YSp7PDsyuhQ4CAug6xkYAiBJQTtWpkiKlKLub6NVPEoy1mpjDZIIiFChqfpYNZuKDCMDFIwRrvwJoUNbYNiwhZ/JEmETSnvMhxlFEF5jbPPsBUqb1BoJ+UThsL7El23zGgUSonlGMqGvAsjRyUqXzeY9cIh4HLLAJF1srsQqp4gNGQRYLa8ClcaLn5GbpzcQHjPgqjI/4vSG7nxjIm9+h0UU7RiyGIErrS0Q/wIxzRVD44EChlDa8M911cHH+Z2zkMsVmBYIxXyNK6nXOFK24V7t0/R6OykLaXBDlYGKhP2J6XyWJfT2YXr8FXPxFXf/Grs3383HvzHT+BL7/0TtGNX4ppveyFs5wCOXHklLnj29Tj0hAuxc9aET//SL2F3d8J5L30lLnnhjZhP3YWPve030c46hstf/+0499KGB286F0/61tfgyIVH8MinPokvv+89OPGlB3Hxa1+PeWfCoYsuxfHrn47znvFkPH7XA2jnTDj+/BfiwhueidP33omH/vEfce97Po/5vOtw9Tc8A9Ohozj61Cfj+HVX4fAlF2P58j3Yb0cw7W5w3le9Cpe85HnAfZ/Fzb/2e5iOn48r3/gdOHr0JB74u/NxztVH8PA/fS7POwvqAkKtqFwyhQIBkTKG9IbCA6YhSlPCfzugXhdrNonu6Wluy28oruT/MLsTIkcDoU5pLkLadEaYteS6TQCJ6oXkeUPhqac8ag1RO2Vw9pBBflbrVLZG83ciLOm9DZ+tUgOFM+LctEGxbo8uiAxbFqtppb5guujCZ/5ks+OHEndwMsb6moi3DkDYhvuKrI/XJe5nxGDDJWzibZQmGlzRNdF81VmIPp2AVF+yzwQyJp8y9mtW/QIE6ii2V1pQh5WYjNbC9FfLBiCV8YGrEEwZGgpfIugYYvg6dI2Wy0rdAXDUn4uqDGyDobFmYkbrHh79xEdx300fxcl770ffXXD+y78aZ192AY5efTV2DjScvONWPPDJe3DoyB4euv1RXP66b8OR48CJL+9i985PYnc9iiu/7RuxOTChnzyJY898FvZu+yjueMe78dCnb8XeIyfQzroAT/qmV2Nz9GwcfdITsD76EL74l3+Ko898GQ6fdxjWT+OuP/h93PfBj+PUfQ9i3eu4+DVfjyMXHMexa6/BNC04fc8XcPe7/xT3feSTOPuGF+LYVU9CWx7D6UcdJz/zcawHLsRVr/s6TLOhnzyFs5/zbOx94VY8ds99KS+VvepQcyIJupRy4ju9D5dIqWLVnAyKnBY/wx9+via5MezqRYBTMaWemd/tOquMy3gXxLhEWeuR3+AqbEN6xFm8RY9JjWkkt5G5CmaqGiRpbVWqwL1xJMYx0Wsx4WQDnia59zPumuTXcq9Z1JmkzBV9fXjXrr/+f3hwmp54TmcpshqKjLM8FErowWNvRH1uLJIB5A2Ua7+up1DVmAV+lQUnXdtQbE/Gh72rbdpUWEVqvDWfm0w+BMFrWU7neERN3xbLTYceJegHqZVD6JThKKTYoIlqSVzJZsMFAoeLSuJMNsJVlqL6XAosnSa5zsjP5sQwjwOsupMQ2PnYuTh45DBO338/+uIAVpz9km/A5S+6GsuJk/jSe/8MD3zqblz9Az+AzfIovO/ji3/65zi9HsH5z3giHv7YR/H4vQ/CbJMNjdEmHLzwfPipE9h95FG4B7J+6IJL4LuPYTmxBzENRXDbnH0u5h1g76HH0BdlxQC3Cee/4Absfu4WPHbfSTz1R38AduIR+N7juOsP/wh+1qU499pL8NBHP4KT9z2K6uNZFn4ESMOT3GP1MAWXF3lmn8+V7NQKRUp+04BgzG7sQoSn8lrqDFQlGyz8mTLIwdrTDpmP0xnyKxwgwg4pKK1X8iu5Hd8z3tXYLDlKLFo7gHU9RdncbkA1vo+eHYV3+ynv2x4z0kOudglzPldlBSm/vqJKPeKdluXOh+36Z3znA9YuPTfisXJb1r6b1lrhhzZ7VWNR1uMn/pDAkkralVsGFr44aJl1mN33h5oC9rIgS03sMpWBFzBHwIgxroqVkpWmlG6+9IpOy6DZlPr5xBxygyvkkbAmqMcYt/sy1BgsKcTJZOQFl1JtbZNds0cFowvQ+z6cwq42bRlWQeGNWLV1Tp19HnfOvgiHzjuEx++8C3u7JzC1gzhw6aXY2XQ8duddUNEXoDqHaahBQVqt+HtxJtTPZGX8XYBsAHi0vmKv8jlmE5b1JKZ2AA7H4SddhbmfwuN3fymVcWYnFMJJ/E0M4Pie6CQ/kWptUCPl7uFpTvMh9HUXa99FMTrDWIUijD6kapPntPijbCdGpLPnOWfxF8Pi3qOVQrNNtucznsFYE+PsVVId4CiXPGuFVQoVhNnAPen7URK/SUPW1RMTwmYsZX/M0GktAqLbIDeAsfo21jxNB7Gup+u++siwHeU3Ro/u7d/y0OyIfhTuBm/0CvT/jKP64JKJQ1EZj3B1WtvEhcxLTNctAdJiBgZ4hLwoUjJyQYumux88DXc0lxAB2ZLMtWWiZs+oNnlgSnTl9zuyMS+Ym2bhjzgOK7Xx1HaiLsNVQVoDd2MV4tMXUSeQZx3IGb05ffSkBCrV7xPYcu1Cy4sULm7tXUNcAKU5DRP2H74f+w+X4gQcu3d/AbswxJBlNWShRVkX+NQYaop3opNnOzqRjrxnubUpPKJwh0DupHLPM3fL4rlTd9wexYO9QyMf8nK6hB5UDmtdYoLHndiOcRJXXtK+oA2xdtdnbBAAACAASURBVCgDsXB1yYHwMuTak0fCzE6GJxgK+LpHbczAOZFVBi20CFkRxVBhphyIiDWkaT12M8RPXoHle0rRhG89BS8ovY8FGjJdPxefk2zm+qXQMKODc3AGY0YLHvKbpD3LNVV2rg3yK5mcMBvcdHFytihjRsU1yAcihR/wLa1aWnREdwdikqsGgTllAEC4dt6FZmzPUogMQ+EG8ZcGVcLWJkgReFx4+pDqCJTCpMsNvVIpqayuhWNVTr3N+a4AoIa52jwJn2oXpOml8LwnPIRk3lF44Cy/h9e+5WQrxaOIEnkP69hlhW3IWg04EixmgM6TulALDCa/X16aKYXd0VFMV0dPkC7Ctnp274vktAyG9xwE1b2S30BwYzrDMzFCFfZl7AxxZXo2ytG54YyrEWD1Cg2uzkYzYMaC3hBMZ1JtCNQ+IdatJfbsxs5Tp0NJUFJeh6sjXPyd893kRYTXwa5hynCgFJNA/ZCdOT0IKZtOqncYrVKOkYnbDw9twBZ0V3JsKMPVnnVRHSv5F1Lgdf+YuuU+bN1PyOOR/OnZAHqDiAYuC5kzEUbrmZtLC4nyOpR+ipdQ/KV0YIFCJWWy6JEujENRvNf43zPBJz1LJb7VTUtp0bDB498Fjm7WMFl04qou3VNY/kyNGqqXJrU7vZfgYKjsfKQYy8LIcxoQahc9mPd0+C64mI6il9ee1nr4b7dhz4bQ0EX3pZX34TBRHJLJNvm+7h6/79XSrwA65DNlEeNaTmlxsqLVLQHmZjP3XNWgO3lhw6sTGM5n957CN9kG6jKmd4E8RmGGal+QAitFX2uteh1LCrNRfgRoJiCestfzbARWZ9Gd+yDrtS5xJDL0ze+RJ8ACMkzBiZEsKsyir6DaDhnRNnxuGlK4Ctujf8WGHsA67BG5D1qHUxEpWyOZy16vpKqn2i3wPj0hyq0USsovRvkNwtwMdBtR+4nAT0/r3diSjtZzsPLZTg9gXMnaCtTly1LsBExVfOWl6T3qNErLeT7LUexBoAQm+j8yHQpZ8iLDwFh30VoJnVxOqIpQa6yioXqWXF5asTh2hk6RDQoKT21ueEYtf689FBJehyMLx2wPvQt1/gY8i/c0BtJ4SZOdahJ84TjKFHQYmPoFti0sY1FdTimuIB85mxtxb7tH4ZWLxYp8Tlh1Y0FYDKTeSh36imaHEksA16HK5sx+GAlnrB7Oqg8p4x6krEy5e/EDIntVvS6VjZqMow8TrJTS0Ms6MykAXBwFbHkzGP9bRgCWf2cK3fmZwJ/Y8YzeZDNWhQ5noOpjXUV5DzoLcXXk5wGxt/K0wdBbeJzoC0ktANnLMKz0KMHPahC5ZNuskS5CY2FAld6T5ZPPiLefgealfZD19NNwea21rFRzHojwCcXX2s7ohRCbEmkXY2izF/aHdfhOTS+8AKZLxayGMhOYsKYyK9CpM22aIKSYdgobRIntlb+XlaxeElRYppZyKz2qJQUsXDdeQpJXvC/osLxIid4TIY/LoDJlYSRiGfKZANwNZlSEStn2CsVGFDyAPdV3tMKRDPDBBZXlLRczyuBDyYipKk+jvAqBxHrviXF3KBSl1BmOshN4CFO0XISBeArg6lqmC5aha0dxKYjFWBSIxTv3/KlwemWR2asDDmDC6ntkrkac70kDtwT4sjQbUnIOYSQCmnXxDOqIVryC9Na4orXHDA/9bCp8XUJEsVgYsD3Kd7zHmjIhkFiVvKQn2EAdp4JynrmbEgc8N7DFXjDFKF6VTlY2RueqEoDg+4SH5H0ffSlOEqiMyhMvQxdrDo9+hphbVBZyrbuT1sxaB+Sh9zhSpjDDcrOuA0pjjhRfplcH1074QV4QBMW1p4VnGqzvZ3wMYR6t8JF4NkvpWzDwxJeQ+xcumeLaKS9DrLFYoGLdgZcjcIGeB1yfn9DaAaiORgV0IahRxKOQQJZWAGlTui4ta7D0IiOkOSRteDaGS0IfQuGXenemMgpLlUox05FzAmShRMLFhfeIlynoY7waGZ+hspKC72A9kGJo38ayMl3pGDyBPlxgnndiTSHUK8dOGo1RWNI1z7GULlAFacjz1y+jrLrkwhq9B11EesbyCQTm8dIri6aGzoXXDWXo6/5wsSssdV9CfuWpipiVCpMeRpuCk8R7Eb1MG0Fo/lyccCrwps5hRmASRoCTIYTOPdO3hsl20nBlvYyzHWDbIQBtcN+HoAEVrIW8MkJQuLYY5tx3CXmJZQocpOm9h3zIq0tLJZBMeWRtpASXu8Vnp+gbB6JIw6e7aFtPycNSt2gJhjsEGiXaLW/IuOFToe8CNLO6kx6AQo30ODI9WMgwMCg3PrvmewzcfvjAGq33VirLXZWktTct9z2UcLrNAIokE/uQilSWZmAfyvOaOPinLq7nvuvnGi9F1SSouY1SzwIEiT9h3AuudUgVw7Y7NGV4RMs1Vqtaep9qQVdp8K0z95I/7WGBscJ7GiDFgBDOuLBSBApLac2twtgRdM61jL8S8hBG1av1nGSobxuEAsDBLvTI84tz416B8ofyCJNoCOQzizdBxWSFy8HKo679c6gOqJReeBby4M8sAAXvk7KLfd0bFCmVGjpmQ7PoXDwj5y7wcijmkqaRII/uqg9fJo8hXTVucu/7yZ3v1nPx6IHej1Owylov1PbBQRA/IAS3BGgbH3EYZmicfTDP9njQ/DPFbS6qbmhQIdri7Kt/pMg+IegdmIC+7scsCQFCcnPDLQpvhgVmgc9YXqoKH8RPifdWMVO8c5TWyx3Ndv6ZvvSsko0H8FDptdUk9AWAuCY+nC2w+j6BUmIS1uCrQqqeGJSjw4RdZD/HoUKW3pQPIyxjfRre1IaqSKQhSHRffw7uI5yl2ON80Phu97ErdlVSjoOK+aA4+9GLVCjLPdOIwOHLI93o1XvW3ck32Mt37rbHR0TGIvZ6BhCGI7y4vVxLhtwJ0o8mBMjfUCk1bNB9L36uL3ALAl9541Hc1dO7Ybg6FG/6sH9ApfDDQ4wCPZsG7ATCLULmRZBM75dSPLt3b+m+isdApFSbvEVVDZblOKcU0uLpHXq6ybI+jbMh00V2+iItshaZghwUlEAeDWzNfDdkzxULO8NounWyzqlRN4OCU3ozTyg3dF138zDhZb8q9o94XWzVYI32PHpdeBOFmAeQ6Utq9yLZxP/0+0iLFdCXnptcYr2r4sm+QE5pIemFRRgcZjV6Ab5WKzyEezqGM80CH8pMglVmyDm/s4ZWO72Jsv6eVpUT5zO959Cgm7ScydZcc90A0Idwrfg2hWPoZ5KzMmQIVMkZmQpP9zzlWU+yOfqaiHsAz14anqB0tBKMfwfXJ5+fQG14cUgeRnBJ5LqnUYR+L490Tc8tpKwnpbtDxm3En9hT1MUROSPLiPCKlrUYy+P7xoiBoSM572jgH0WmhFfZRMqc5BcT2G1kBdhAA72zrWFPN8XX4EXIrYkN3eMXK0QpLMKxorUghCDpyz35/Jk3dgsrKg9LG8mL10lIicKdkfNQGfNtj4f9FHtnMZgwiT5sEnKzkq2Yrl8RaxwSQmY4uCY0VZoy3ZupSBZDScWYak3Ut7SayqbCRK1FF6av7CKVHpbWYPWe2ViVKbOB4BXdtIv37y7uDNOPvecl6useNJXbvMWEKwccQaEOavNeuduqpOQlcPcE4DJrQnfcHCzYksurfZT8OOW5c3+KWpxYV1/SO/BBzkDXOADyjsDLWhqXBIYpvx1lISMq26MeL5q5AO7uK1p3gGXfowfEIBZKV8oDUzgn8TRYerTpoVqFMlsV0DR4nvIj3EtnWtygAqQlv4HXKQRRWlrnk9krkhJ73x8SF8i7q89ng26IRxOhkcGw+mpUFhQsLLlx4JeNoGH3sqJwkkusLke5lMZmLRT2HvF971YaNTX1ijVxA1nt4MajL6SB7MMZCiltONZtZEzb1+oCvhIJthneLIUBNnQEGrSzsg9AZYSAlZdPngg9H+fMTKCsvLPXBK1LXqq+hEuJFZohG3+md8WwlgVO1N18u9BHFyA0fyg5TU1T6wDxDOISC7RcaxCw2VDX0wfhE16j7wTUOCjWGyFLt/EyIy9x9rWkgvO+H9PEIHBc4UtgW9UhK7y81UayXKWqR8o75Omimuj0vhsXsHfA9nJP42e9sBabcs9zLewtEaBtK6XC73MPUtlE8F+uvjXjuMNG/GONNGUT/Fdp4WCE8uwGlqRBmTFPrADcRyRGwsYzNsGxZHjhJq+CdyBDw56KLpmqECZHBS6SZV/REY2R1LQZFqlwvacrA7Puwy14QrPDPS7eNLixnRpdQKFlXJ7AkgmekcWWS2Tp7rgsAb0G/m0qohh1F4JQXP3QkdVBSu4kqLQGYU2ro3V0NLDXBbM0OiIA6erm+rCgEHzlzQ3pidCVT8FtU3Z9yu8nViIPyA25jzWBXjUVxHRkfeVupoCvmRXJGJX7bamw9zHZgbIOsjyqs/AVI0svAOAIF7IWJD1CXR6rEHGMVa2h9/AAmnHytkfz2s70soBOnYv6sDY24lEIgSHzULgQFQocI7goD6IAVWe4w9Ap5VBDr5htU50KDV/1I0Duud69QqSW1lXxu7KAFd4o/FRoaKkcJDUtwf0xdOXuEgMQriK+j3p0KJx2GmaNp0jvM72AuqNAKa34SE9Zr2mBzFhB3uzAfoYMZHklI7eqIoAiE7ZC4stlqhJcHjR/qxhbtNcEjIBQAHQzNSoQ8gTC90t3TQLgAgNRXYLGtTTbYGLbcwkygOp4rJhUXglqApkUUPAAply7LoOamG6h4ZkBEoothWMZg4op2IaDGwuJWlKxQ4Qa29mPTDppef3s9j5SSVOgleNWXUF9vlZtFAzvK+bpIFrbJINVn80Lb5sSbOEqPN8mJaOLSSWo2ZpR48BW9ynAaiKMwdXvEIvQhj+vPZq2lPhYvi1vQ3KgWh8JvW3JCNmT+bSiipeyl8yW/FTpgAy5lzy7qoJF/mIXMikkrdpLfrfXj5TnqW1IY7dS6tBei/3sebfU1Fd72myDHM7F/6WXI5A5L7+Ucd2nVMhM0RfQ2nLNLWUw9lJG2/gnkl9rE2b3XhueVtZTCDW2MC83l6NMQss053Y5e2i+PcCHrkcZL9HlpTU0GNvbDSGFd2gIitY1CoIatI4HBCDLv1W115pDGLpiMgybDvds1JsxopXbFt/ToCnxJme2M5uSTVzj/gQTVfHpkpddz42HcI6kOTwtYU/lVfHqmmvtRMfR5q33BlH/9ATWvQibKJQAGZIZZ2Nr+nc2NPIFK9mHoAXUrCGl9gAWBgL5rAK55SnJIxBugOGZ69allLchBH5MP8uVTnZxXvpym+udFHtXYV8aOa5NCkHykxpyuIahj3XpaPR0CU2KRTiCp/wmpwcyRkueUXotVrKfSs09K2pBI9oZ8iXgLq8UDJNd5fPC6Tocqs6OWqq6V+WNqahTr927amEEcFaYpCghPbEeZzdro1KLwjIOkktVoYUApHDPneQhudSyxKJMw+fMhgT3gKnPIeNQ1tMg72T1aOJhjQokv1sKJdbXbJNxZlnsoR2byaIXMKZNwXCQGau5yn2RmraTLG8iINGrCuHgbE7uVJNEJfgkd5pMRPVKhKxP/NNBmjIEzg3kNKu0cmQnIpxqEGZU1qlo6eFGd99LC9atKitTcNM9bfl+VZptueb0OqRLMFGfUDr0PAvvLkubBbQxnFCaVcojhx3lkOIYSVghThH84ryD/dtd1phKPD0jEdsYIPAsQn5bfren0hqKvSAzxf+ySBy1tlPpyDYnLwRURvL0pGDSK8Ymb1BlGysUA+LZAr5jLawm5bjHSeMznWBwekde8suf7lRQkx2gjM2ohkEypmVwlfkCdN0FiFJ+abQiybCB2eRz74v1fjq/MPPkRHkFXkp49UtpH6VX8vbTXc7P0vK4L1jpcYzWopMW3azGvbtzcF+29ur0YKqNn9MlFYW6mWJ6bYZHk5Om5iELVCRVoKQuZRwTEmMguSqFfSL3YaYGX9BLspD9NRJsUgPaomGHImC37TElytoXpSxLmMZ41umNxXf4YLV99EZ6zz0z5taXfirJOMvQoVyWqmanOrkhEQd3gpHdV9h0uOJZPyMMzTSyYv+9aMSyTljWU3SjqyFz1FFotMCmhJlexdp3aw+MGTXG4MkskEIll2Dtp+G+oCtkQbExQ5mpxJseH724ugzlrQXOU7U26jWS38vMlsYBrCpjaExZdkCYRMkGM9bkiohR6b5fRopcHl36ZsC67sEmra1aJRToXWS7UiorZSu8kFiH3s3SA1ldHiG2n2fIfZKHxlobm6e24+YH2ERUeWX1dTiYi9TGphVPFBV52N2jjLkKjuLEzSas62nG0VX1mD8jd3nMvdsEMw0VDpB0EjnK1/RSpM2zwcwAJrlFReTcdrCuBHfSYrUUhmR20nrDldqKPwVjdafGphyjAMAlrX6MBuDllhLhgSj2HKsmcxiuLO7onoMdm0FL0Pf5OdHO+f5Mz8aiOr2JmJU6DUSgLGse9jgJcdpLNjNKPEZeXrcqlpJ3pueoWA89wc5mG8wThr2mUFI+6ns3+b7xi/Uj7lh9D1Ojos7GTBF6dIZ4MwcYj1R7GaPW5MlYkeSspeyaNTSftmQBsOqChcJxOmuMWpvRfM41ty5OCPckrXkohjZtsiRADXE0/jLeFolNuA9t8axlfc5kB7D6HlP3Vnu6FVpFbU56HgNuUdij7mThNxnKkW0aYwc82/7Fue3D0W0OK7sC2VMiLEtaRn6BmpzWg+UVKBRZh8W07BYUikpUa2k+al+vNJkErzIAQmNXRCPyKa1mXFYd4HatiFxT9wo14qJu6bbhNwUoVriiy6DcOv1cr0sl4c9YdzwEk0fhlB+1cBupxQSfkOokzmH8Hkc0oc1YFwmCBScAgyu6pgejqlDF/4l4m0YUiOSzog+t5euyKnNAXkTXLBWh70q1Wr0nnJkSYUH8B2XlYw/CUxjbH5jHE+szu+Wt5fPVl3NE+svL8sG9L49nTaWw8sJW6nj0XLlng8KW/ApPMspDjtRks+X6GQzr0x9JfoktqGMVw9ns98E+E2Uw6Ikqa4Iucdj6DKxBg7UBKSzdH/C/eYaUsQZhgAOQPJRX6Pc2KCJ5vHPEvzOUZmokeUT1ZWecCUzMjUfONxaa7ey6yqDpTiqeZL5WaUUofhYpBz0FJ6ncEoBWaTbhWaFJkRus9JSoyWODlgQJe4fZMMDGVzTbQbLgvCohUxDT0hUOIiJRAWelIqq7E1BaW4CmsdtXx2SbJCplxskGpN9mdD8NzZiMDAc9NSnQbAAz8fDD8nbxMCD8AUiCHM+wa/6GC5cYlWOFcDEGAiXoUGEhGx1RAWkyXPc9aOwCXF7XzMyFBJRKUXM+ea1lQKoPBGN7eXviKwDYwraU6bEZDZv0hPgC0CwNtT+ckvLuUNf6YPYuGLuAZYGk4vvBK4owtMFdU9elND09Tgw4jS6sExeLUHYq2XSBnMS3eke17GM6n+X0MsbeqjBPRXON3mkU/yljU+vepsJXaJHfI4MikURxpwY80OcYSrMbJCDyHiruP6OwZhCSdd0GypptsBJQy08LG7AN1r679QzFocJG1NZOHs266jM9fnY6mIchzybco7iYmhjljZaocWhwZmq52e5Y/fQQKhnW9VS2+JcF7lgGJQEkZpBdysPKLxx67OiYGLd6aLA4DGu0jlWoJqsuen1aWlofb42ga7EHwXOZ20F2oaK1NlnE8DiW9XQIFMNKhYbpUkJt4JmntxjDKBxI+EN1TeM+oHOtGscXLfL07lIu3fYCd1gj9MSW11KKoX5JUa7MVpWLPwK4yjqoMXOzDbrFuqvfpvGyCgeZA7dCyzVCJ5RWndksq1EUkmtZfnm53SZY3wbLM0SyIrZFNkRh6hIKoMWwq5XlCMb91+S83vcDP5HXpLCpTTAabmVTAiehV+6OFczm9QUr4g7lwDAPdrayIxWChRJYt/ZnkilIrw2ZGnfM1hpaZyzLg21WVlYxXoFOcdknxqlucnkMm3aYF1Op0aJES8sLNVdZdnPx1jdQx+EgIYmu3TBPrf6utfzzQriJd9hIGNOQIfZNyFUqVhOoGdpY3bkCeBpSyC4h74MQr7Soa1lIt3Rdk1CGjpZpvnI/Ic1uccWFdCe11+V1IdcaHiAgUJLJPQrkSvyiOljlpHWoG9kAnKYVrYsRym+GUsGNKbiGGWrAk2EMzz3rQtzy+TEcivU4bQzxuE+2GULDwaoBmCeB3PGrARkSGcu0zSY26emY2auy+l6wZAEa4lPMYoG8+j4XfoTCLLBFDCP/wNTsd83+oTAVVk4w9pBtbWy6U1kcs6HK2TuxgFBKYpvEfrMTGRqJfdOAQcjaM6TNcLYh+qHI+ntiIbnnlKXyBFnnkh5QhSCFUcQ7hPyyd4YBMzo8hKfywcOOQfhFaNFlcFNi47NgDJE2CwvacsPlziuFJ2ETcURkEb2e2RzXNz0VItle/SaEG4w1/UrnjekkCVD1kZiSjBKfiUYqQvIn20GW8oJgmkX60PWstoGva7avWyG+yUyMxqjQBneUlPhmc1jDFBASZKCipRjRJ4BPgLC8HIUjk21If2cWyfZTyai1W7OijEvgh4NNxaVwpHAKcgL4Obfoj7n2oUGOlDvOOPs4QDTbcI19eObIhhwBNuQaxrhaVnqL40ALmZkYehJVf6KQDYBo/2gFJo68D4YcOUpyBGHpNRjPPh6UJAPKN+fdNM2z4d/bsAbiCvJeKhRS34lifTbul8nA8vurnUIRBEejIBAYYMMiU18QtStQ7UiAyqk85XmiQqy5HYxwlvdKRMJmDb1NAeuK2y/XvLpgibLMPLVvAzixuQsXE6kgHWuSQJju7H0PnZegUyhisWWdi8e+oLvK0xe+3BDWuOpWltTSzTxi52GjunP6talIiCPka/WZOgNAEo6j234KTPcFk+1QumIMY/f9AVmXlh5c+Kx1UQpajXk73y2whE4lWlOzexDZePnEkygarqLgwAi676H1vfwOcJ8jxTdlOGmI+pRwy/dT+YeC2oGowvFnniGFCtDi9wtWYTr0ms6sFQLTyuHaCn9SG3rLZ5150SvDReDRqlYoL12i/BjSt/Fsz5Co+DLxwQYDa12gUFBgNUMGCICkBklZ5tQ9A7JKmOl9PaNjqWa9UE1IFQCWpQ4a/IolQ6DJdjJ9GdY+vG1YT/kZs4/qDIdBmUm+VDfVfR+muhklFQYQPJ/bd4emTfS0sESAOZypIOaQpcVmy9lMlbGdhzkR20DHGWnAkU+hi9WqG1RYFAJf1uO5xmpFXiyNUTPbIDv9MD88ebUxy3ZsslAwuK1wV6q0waAhSSEEk7OrVIvYu/mMqR2AAVh5aTzTVh3rkJbS+ta+HyAZMwGRymW2SJtrdYkMhmbxHd3ZIRyGqglZ+X1h1Vqb0LvQ7ClhsRA6knNoXWItm1QwDQeHoTMUIF/QbGdIcxYQC3d4mwchET9CDYKqFiW8uohXJ5vjT0naCz7EaSjLo+pggwEtlP6EOTghaZGLCj7WaUQmROGhQbNGQTBbXcHl8WS/Eoh85lhdZf0iRW3SWwjXnPNaQOPmpFtnGn9K2U7iIGU6iH0WdjbL7Ctk1MjPSF3HfrQmvGXOd02QOn/fYEnWkXckjyyaFzVXKKSmQj1D+e7V91NKfe3hvVTSoCUmqDLzqe1ggWgIZCEbSZUwCDpI+ZAsWhODc2QBlt6sg13Teys6eKXkKq5SiCINred5aXUBeb4SIVY9wF5tZld8bLlJJnAQ6sTU6JkEYSs0MT2OvpsWuZH4o+nnCWhpZX1l1aOsVSe3wdOND2KQ0l/xLLX3i32qFJOowCPFPF3cLs9mSOd2zfOYhn3tvIT7mORN9P1ci6dyqnSc9hoCr7ynMOiZCpMqJKF31xfm9+W5rWkIbDiDPAvJgPmQTiXO4jIgBsXWTICSK8IKXBqiVCd2RhrSVfpO9aTcd0liWvStwry0ivHuzVoA3Xn9J4gIV3E+MyDu0d5Od4EZJclsnU+lZDuLB2PA+5oXO7MZan6THpmA3KErFrGECFuiMY9GcoAKrlNG5BEYPSqH00PRWe7nHgkU7QMjO+jkC5wymOneAchVZbbRO+XwejS9jH4pfgVUqUcBhEhNUhhnhiPFacCQllERF29LCc+Aviewlz+jyjlZRQq4qWvPlH9nemkJpsql+ffykBLfyMtQLEHFh9KuYeGn3ItGTKOZ4j6CeW2H1mPOdQsUU/pTcacyPkL7s4DP2hBn+tYeRB9Fxc8FUlb0jLTuFfNX1aEui75fCjZj73x2Q+IfgaJluDB+F9zzOWkaElSMnysvtJcsDHyIctnVKMbzny0WYgiKVprud3EZwlj1Psovz9GEkwk7wraStDJocUmphLLSsuc5jBhXKkEAmebHWtURaXjHkEdvIICcyi19LoVrynhV6KFNGPdU66hGUL51z4ozQ8wj5dVS/vL3nJKWZR4ILzxIYlVU2HgH5t4XM+/UvitBPl5iK1cuPYSB/FPuZN46yGpXvBzuW+8Lugpe8md06NHuLjZiTWq1eBQKhWK4i6xaudZGja2zUXYgSn130hLEV4p6PSC/LN11ElykgMLCdRAwARr7dPRYbzRRqaxRfp6CobhcQtBsk9/hHg1istcGxCnwvGiZeUguBCAOivHdvZXlaoiUWV44R6X2PAQ29rZCJnPFt+KuqFw59meVl+eRltbZLetuzC5TGpyWv/tCpul2psMsGKUQTpFhLsvu2wFSq4s9e+Ylj5R2H6zrXhqKvjoEIhtYeKeUcOeewmFYBz4JktZe56Vu7uqk3WjRY8BUZUcAY6VdrL9c97E369hQuCfHZvDO8k0DW2kwLH0/yG19QXX0Iq5iPeVe93RUcmPrxW0qPSJDRn4G2hwdy3V701vpqZS0Nu+Obgvm1jZuqyzCBuqqinQtwwAAIABJREFUU8QScQEG18bE/GKL/0SSR/KL5QFn5mOLMFIuaFUshhKIydLOoqmyQuV1gBstDR7YR2VVSKgJTzkVUsX2BRBpU3NgM/ESrSc2kPHuWjMuLUEznOHKKeMzUTH1rPKsdngFtFkf3dva57Sosh5W68kxeA6GNh7dzYb3QRa9dVE+Yvc0ys+qKM+23mOFo1ixIlald8afnWwcBjXl/ssr00gFgebxXZvI7KQ8tHq/RPoxyJMWzh4l/CYxFRs2gDk0PjG9U6aqm+LvmpyzpdxH8pyUYGICkqQEgNmaAMoU6ZFjVkcypXA81iKyYL6jA0Jqiv/i2Ue2UX5r4BSVPkq+6i4LwI2vTgM+LDJBS0PKUK7XZTx7tqRxnkeurXXAzGZfV9Mhr8nSk8X11GDFdMQgWHtQjG90rZICzi+tAyrhNzOo1fwgxoPyQP55XpBBIYUVngfrVHGsvqfZjBUcOGwb5SaQFtXUOGXoD8E4PHkWqQRmiDqrvpuOuJCdBBzAM/Uqtl1abJGuGAvGM3Usg9I0ZZQAwzy8z7iHowsc35lr5juo0hcZy+sZ8vaEpPd0N2XF6yIbyT1g6pS9ITNVrXBne33G9SndF0SjNnzX8HlhAqmcCiiO9dFKsh2jWVlDGZBEh7wzs1bM2w7haTrTGqIUPyvF7tAA5qpVqvs2ZghKzoYqTT4z39HrU5Klkl+Bs8FpSTAdWyYMQXIkQ9PmAYKlEmuqOeHsW8j7KAzNMYbktZaueSTAlvyOQ5+ju5vnz7t3nwWuuK+YZDkGKw2jYjalApf8fAJPUEy6oIEXRn+W2lYxrFDpYId1jgLQC3WPtA4s2G6TKhMT+VVhzy5fSq4YC494YaMcdx/dVmCgewsFFsFIFYRVmKNUmmJ5R/Ba1wRSB4nHqCQgxZb5aQlNXcIO1RoMBWlpGsrL0EUalWe4z2NaWFdlFLU+ALzscG5jPQjJOa7zrNoHdTbrFNLuBM98+9xBlD2WyUug1ngeoGvHXqZ865oxJSkDpDULsNaJJr1bISbSQAlHk6KyzB/RIg/P1JBnQN4GlTyfVciAwPcVhk2epVrbieoPrAMgzzICDfam3ly90pJKmUboWdmQ6EHSoTkskTINXpG1A3lvoi2fsn5VWi6vzxlSqbpWf5Y9VgYQNZRB7ZV5hGoA8o4Rtchzkf9vDrQ2xW6GOxJaQVRgEapahiFIK0EkImNPOAucCIy4q9y9av3dZqbgVOy1EDwRuDZXbtiwBeg1goAiowSOYAODkqSoLXKRJalJab1w8SZanNEV5WWydUsYja5s/Bm3L903Ak9uUL/NyMuLPCN9wks0hhFQX4qho9HW/1T3oWR27Ed1N+K8Dg39gdf+8eerQ/aUz8gKz8QXRL3uqTydoJ4KB5sdxNR2mGreQGlig/gp5RmNWSHN8AzlwktthubzMCpC1lKh3/BvK1deAmi5nzwXCPugjHEdmjDeKMfyiIJo1KiIUaXykmnSAbKTt1TckLa3BMoZcpH0JDAVQBT/AYTVDGiUX2UYKHvhMMU5TW0H1msuquR3m5QVe9OBxMgmKQoTb2Zi2NkpP1Pus0JY8yDbCZvyLAlQKQOp5Hl+cX/mvu43rLsIFqGzVF2gzIQF1VNi/FVzJYgFtJ2YLGXV8t14cToteJf18G0B00EmfdmXmCWpdJF3BP0YnDHpAKslK63rbPy7UFseYKgTAte7iqIEYCp2U8Mbpv0g14vxLy91eQ6iSo84DCjMQxMZYST8vQ2UXFNfRFkoYjPmpYThnrUyku6V9RrewmWXalFIAjcWSU0BVHnS3/LCxVpIaINCQY0jYEig8IDrXPpuWCzNCg2YEQrFqu6ASqsvYWGh0AKoilICkl5zNpzrlDGR8lvYPiB4H+K7LLzQ4TE6eoQmDfFdNmPBacqow7GXa5PFrJThytBbtUmqjpX8qnCsGiOZCSAdSYsObxWidyz53wpvWnZR74NnxAwjOsCUvJToxKlx6XFrBggVL1gMp3V2DSb34J/kzBTKe5c8qkCPtWCVvUEqNOS3OsZh4nNrs4cbggE1LxBSgE5RcI2HSc3PmgdVmopk5YznGxubhutfM1LlTvNpFIQ9iOIbyDerYIlUF7C3HVTqZSYTAUruuhDuGPicI/kGAM1QvABDKYM4mClwj2zAMikyS9ecD6p/k8W4jXrL/tbl0QFNbQer70KoNgCoE3d8Vr1E9or45IDcV6XMMhPCdQcGNQ6+WTKers5USkcyNEmOwIRGhbBFUhMAZxu4msU6YGwKZK6aHa0pZEepOlHX0yslYxcW5zwCrvEcUe29po3n31l6TzmvxIbQLj2N+pkKt8TfaJgwp/ehPwEcnXIm8l034WSDB0TFi9aS+KRJaiG3a641weAsI6+Vqn6pakjULMggL1bzhRMkNaXBhXmMoGe9d4SUA7jv8b0Ozxomga0jFyoBdQLUcI8enCE05XZ5r7RTsekiHhoBJI3T00uDmZLiPUR1otxR0amBIBlF+bCovoal70KVjmBHqG4q8Z1CeL0ATVmHuBg1Z6T7Ong6wTFY2DYetBbCBsrDURqtuADrEHOn5+OaFRFKcpWC4xaoWjNTWT5MwgaGGBIwCzc4sxAjiOkC6fYB30dV6qrfY51J0Lt7upRBzFnCagqrgNPaGM9TaemV/81zRQ/llbjTkvvlDBE743hjP1CVXsf7Bh0+2IWaDKcMBmXJKjslHCU08MgVYepXPT7S40shzTVmtsXiM2tnDxQb2JjCK6QMvGOCQgeGc14ebo0bWPJ8ui2pxIOtfBBVUhCh28Syd8mtnSG/zRXGKHwNr7LkN36+WeB3CssVFqaxMct7OaagackAAKsD1c9ihdELiZRsy/sZjwtTWYzPqj6GNfS2BsoWkapcmilBwBF0KuQ3TwvhYUzD75HWvCZXybJNW4fdWBHazIRnsxCmimg61LBFqb5Kndpw1cvyaAWq3hMZaehgnPRzCqL37H+p1ZUr2nOtY9l+TY1vLEsvV3xuB3jJo9hMCL0hcvQd+7VfHv1CmsRHue7U9PxZm6CMR5xFq58fPKXJKhU4WQzRVaiY3cXpxnZeUMXh9UseARWY0ZVGMVFjnmiFpon6w6CaHT1J31d1RwO1GKJ/K+yTN8hiMhaDCfcJercyJ0CNMuAqSMCachasLKlYrWPIKDkc5dcgoFuFghEGCWegx22SNxuwopby2zgoKD4XNSFmkVCO82BoACFua8pvgOAkAfoGGoEwyrIwCk1+HwmH6vaW2Sl5q1TYKqeXVy/MRWFWKKsOmHpv1HvPDZNPqBw1IOCQdQyorsWrGsZYtAgXOm6kbUdIWwekxfY+MPWGS6g5pmm71UMBPZu9VnxZsaxTEOSuBTuuCFxAaOKIy2c0o2XAHtAO5LNiDRH7hiehwp4qWnI40WinPK6oqeeeoKL2brUqouo29DsAAOzm5zsvcLc1LdlkO1sMPjWnNQuvQ6lEuaTx3lWbEWcXg5lExcZgeeI85BnSsvP7AYWVHd3ksk+pMCIPvyLT1U5yT/5yQhzb9OZKJxbJrIxOpebCK2AZui7VwPFI05A/a8jmS+gZJhc/oNGdbnlhwOxBgNYhv/H7ajtQ71SWseatDGlwgAWKImBpXm4AxnmXiHWpUTNSfqPPhTA6tVKXZ772M87PF6yg5zHS5T36bACgR6jarDGTxvDOGjpWrL7L4kgMil20fjaSgmpOljA8bbHZ+2rxwqSB9g51uw6Phgwx0qhzFB6FCbwYE7GFAPgq7kowL8MdpOXK8AUqCtqhZqfG9JZWrMIQxaNyyS2FpdsKUcqMBygCUSgpMJ5EunHqiRGHPMPTEk0lTNiQiKbnTuSWlBdURCdhNiHEE9RTg8QmZTQwzL5ERuJodiCFdZXXk2428iJNVuj/lBahupE1NMy2U25lgqUUe3qKGc8rparPEIsSbtBM5yaPgdT1gYDnVAwWGixkJJvGxqrkRcoLlLExNQJSl6++oOjaxWQV1dmZolXIWzhb/b1R7rIWB5b7qT4m0WyG3bx0EmaJ94zEqC0PDTSKlIOWeFYrgJP3pzAlGhbXfhTHZ8Im2xfwVAF+Xxqb9Mo2yFEANipUNSNSC4G2pVgAyVuQy+L3CsupcG3Kz+letiDg+exYLSw64ETu+7pdxhw4gazvUhqJxVqRLWDdvDnxENJmdbBMW62Zphlxh86NtuQGIC84NTOYV0Y1aNHngQgpcpwiXSo44L6P1QDHPgVRE8KnXFccIOPrtGxMt/mCVd5D1jUo5ajYnx6GMh8UAK1t0u9ZKj6mUyHGJZAXaaQDd9+DgE/1RwgrJsIOlRoW/vk+1ANk9Nrg0UFcLmUCqukFWnIIyjoDyTtBL9CaWYAugFhK1IBVIw9NncmiPwJQma9w6we6d1fVatv2TDPUGcA+yEld0H1KT08BiVnDui7lvoMhqUfCXHG++wojrhXNhIQB0cwos6dQx0VaEoaC3B9RwZ2e51h7pCyM+DWdOFHJCP8+i8Uov7odKZe87HmuI4dC96g6dBV7V5mbNrxLGJWUf5K51jM8zDPlc4bDTTwCQ6QkYQnK6Jdc0uI+cDo6rYub4shoQrMqDeiA+ijEz4niu9Tmq7MSFMezYQwtX82jVCl6XIb4jDALWW8AydQjV8RmrALRHBlCGHPSirUbLyoYQ4eOF9+DFG7+uzgjRTEXviKuRuPhZDqZ3o2nRzKnkhizDs79FmaTCoohoWJ3hWVFBY7sjep7INzQ/3tIfnlDkIDBIZZfNPsJzkFYU/VqJYbRF2IDQPchZc6xlsVncQBqAD0SqeQR0ttID6UspeXfEfCUJ0OFHLiJPApaza7MgEFxOeTB8WwbgoAWlHAxlvl32o/MzggTWLnfym6JG9QG+a30v65wYi6JnTVEWwXQaKrOSp6N5q+G5yGsbVUNi+6cjCVEjlRmsby2+P8C2Mtb2GCiJ97lSVN+0liYwlT2jrWGWRbMkGFTLkq/G12/oIPysIlqN9vkBvau8MUTjbfU5uVFqLQ3XriHZRdKzDi/s7lJlhPTy1GdfmQM4qV6axiH3Y4uriyD+4rWDkADaLcK5AbkPb6jvJ9Qgg0jg1Tf26DCIudBTOGa8pmudWcKqtSvekUq06EqRh11YhdKaXFtSm+FnSaewYU2FIKdzxsuolPYxtLpsEqx+i2r6OIzCBcRThPx9EqfKdYh19vJeyD/w8u1dmYRxGwdBx5VxzSFhEjSmBivSj+qibObvAZ9s1ztqW5NKl+U/EGhlOd7hZ3UjF+jN7skuzZ/lrhYYDmiea+A7+X3l3/i+We6H/CJf6I9p5w03TM1vWEWix3KYj3RW6R3eSCebz16NA6jLSnDX5XFca/E0lVj41QSCa4z7PUK4UTbK48BdEeHGFWpwLgo5b636MqHglFkDbYFPiIwsQ5l8Sw31AjsFLA3xmHhmYQXIICs0milLdtWvBXgoSLyCbAph9Skx5QZBh1kgbJjF+rZNlBvgYxjIQzBKkzhZm4xPiU4CfqJHddhPuWBRTw8p7gn4q/vHHAFeV9wMTbLKiy+wHh2nQIpF1R71uz/L+tskmTJcSPsYERVtTYyk9Za6Qo6hg6kK8xFZ5ZayEym6ZcZhBbwD2C+KbPuepU/EQwSAAGHA1xOL84czpxHj5t6k/bqeqXVKWlqOtoUwY04QhpZmCEaIZQf8f/xr7OgKrT0NqA87nUZ7csEsFMOTiNcMmFPIuvgHvo4MKsDZsOxsCxYj6kRChfOQRNHyrpVX5zG/SV9eKRhveCucIhTypkLZLAa7lx6RIlkZTgec1vM7+yCzjIkT/+7MKDJGjaehT7ZECxh0JFNU+ADg2dDbdxmpZ5VNQlm/HkiM3cVTO3dgCZlzyETlw5SE30vYCji/jmQG+GnMW5QqQic89XK0S5jjmWTr8s1I6duvxU458FAzjnTce+3iw+9u/Nfi9jVStF8h9q+2vJyfXaZyAJ+l45eGCi6ZjdqdigsOj/DBynsOCBaOXUOHOWnYxcK+ArMyW9zfY4RhTwzVbS6Pyt1F6Btu+5hhfyu9zwfQ1kvtigKPfNVg6nrWVk873s/nXVoZuCxFsHcHPcie5T5GoYjMfbzGuZpprpBTUoc5JSbYxJmzWidj7kQmTp/9wQ1eX+IezXmTsEnhLKlMRfD+J05zpZRmbRVMow+AcqGMzITwijNV8qRrY8xe/3a2PVn7AmBbaR5Sp5D7jlraFypvwfmlJIi7rYqdnVxtyv2nxZoQw1+PEZo1iFopxVjz8EsXUhGlZ/ZZJFVCJXxZU/m7anZOg8Hqglz+CL3WnA656OXRm498klgVMpawcns4OZX7vhMh6l3VbFzywVPkgI0vZsEUYA0KbS50FBlw3/3GSDtptdYeh9N528ya24hvmUp2YqrX6NydQqiSBmnIgaeA4QctihhTIjDcXk+1qvDFJ43d+8siVJHzjVTlYnKR8Xm/O5nreMMHK7tIihVWvg165lDZcYQTxraftpBVCuMYDwLu8Nqr6aBx2i5YTOTQ4AyOhQKvpXdzpDXpelYtmsPXUWIyw8fesh3yG8Iopx8X9lzZb30Ib/lCbKpOJuTeHcyGewZ3gN+Sa7Wp9/ld6qla31n4/PnI0SmUa3TarkJP+fIJmeSPMp88l5x5+woZW3aUuZYqe7i3SSprx5EdHrQy9ysz6JgEx+evQDYRbHCBCsI9ZJrVGI8jx210BcH7HaNBR5LXfXJAYzYId/NX9Dszs7ElOs1QNvJ9cnDwq9/GOvuXSdCWvFdgFNCFafoifaBGOZZ5nrPhgJB1m7Py5JemEB6hgH4iM1ztuelIWlBqqnNZ7w1hWn0/WxqLkKlZb/1zj+Fl0AyBuo9soK7K01qc2m8Ef4mRdg8kg7REPTz8B08iQE52ag6dWvwuMPLzbGVYyzgWchGZXpx0MHMocGH/NrT8KQUJnK30kfv3M8xni2o6oTZAObs0ugTyvlZlhDtHZ6e1rUub5wlP4+Vn7HRL2T4FA6XEuDeLSY08kF4eOpde02hSXuz1h3SUki2nXIUAAcpM8gmR1zbwMt4Gidbbw6tASw0iCUfH9eNTN3B24u795Tm8qDVkXpChid/iSrLHhseTT66fZ7Ik5OiguDzHEooXeWF9C4MUDneBGAfCt3dpwycPvtXGbEjo5D51ht6bsp4QXXrzsMLIpUsC03RxXH06GxFIdlLlybHXvP5tPES/JeIft76Thly0tCzdrVG1/oRp3fDo1FKXUew1WQcKVwbU6QfaTaOZ9ehwDWmKdqr+anrdlcqC/0mVRmrT2crP+1lIx79nHiPIP7bzx3CM6wQoQzxu5W1fkZ+pymwbHuPFG5OQyPkLUzdxqtjDMveJOYIbIPM0AlQdvFEOid0cpMy1VWt6dPegl639blng3/d7ltaRhXPkTaKJwEurVHd+9TzmY3NlTf37F/VQ9b3R56e/LNloVLfUubLpQTvuHGssC46XWuMrHA/z/jtdO127z7UL+D68fC4ih0jIqg8qN3QK5YXl7JvwCkOjNWxQ9TDd3mwP9/38JjqDJLXYeRiFL0NYlhQXD2pIbIUkOtDc2UauegiboBWMR4Pac02AxKErXHz5r0RcMNXbeiiMzOPn6n5CL4vHsPCgzi8lpqJe4QrJ8RhmHAq6plL5Rt/6vBl4nvGOgoRfd0P+rfHF8dYOmxUHq33qMmJIwtSaw/vRHlkFeRMiOg9UXOVTQbcgrDUCqUxQh2TizkepihhODrQ4S9z3aG4FS+ZgcG1wNU6k/fx/GnP923f7NjlwVTi6BjmcbX8trEyoA1xDFm1VzGQAZJdXq4Ia+O2XMUxP+e5PGqv5wB088aadugR4ePRjnDEH6eLMINn4laj3DDhKF8BRZcj35NvQHt/zfcIlZSVB9a7gcxytODFuz+F3dly270kXWa+evK8Xv0c496OqzuySLyJEAzK3D+Z2rGNZ0hkKU6SzHzW8w9LzkVvpxAxW2rACgOS5q/8/lzE9INoc50GNINUshXFa4zaIKAT4263NAnn5VcZyWOsihBtCpduu6ppSfnSo18qFN9hY7MgVyuuRAh01qyALdgFDpoAs1GcZK3V92fcZL9Kfq+WTeookJEp/77HrdeZLYBTIp2ngWH0KX3AW+aZwnM1Xnn6+V+9yfHc/K513L25TRB9GPU2JITaU2tT8zzZMDzgQBa87gOuSl05nVls0QbHZ1NGYDv9m4RxSytEFSPIaMXKM/C0q19nZFbHaYNqmkzFx4PleCOF4MpuLlkFk534vsqStXVti8ywzxqRfdwfV7AUBVNwfq8O3RlWZu8vCVU4D4VANKTpuHy4vJrnLJzn6t1zLD6IuQ0iQuJnBpnv69jAKT/vgBLP5wcYrG5T8yzTItChVubMz34f1/ZCNArvVwH3bFDpdVG1O0fVJxgG3+x5vYxFjMfTLfHyzPjI8sCaps56hE8S4BiKTvn1ri4bP3dNhyHahmOJDJV+u0fTvVt+J8M34xzPanQAY3MSywBcz7XZvf5q+R7PBTlGZ8bLGQLZp/y6PuRYs1obGjMPWHziJjrkdzqPHRKW6Kt1BjDzkN8uVPTGak70gDfb7jpxLrxx3PatV09oUaiJ5R3nLrsyjW6Xu/PkW/dRul2DNussH7uQB6pMBqN3Xx3fgfKq+eyCpPJZ6FXK6ANp/f1x/3zmKsh0plIAobPIhD7y61Ve/9PGpqIOd6mGyZc4yKehmSwN83aGdLjX1skZJ70FWESDeU29zrS3Jb9vg324/dMIiOuZQO8T0JZd9+43Ma5WC27LgI1JKffwDCaedwjmc1K2XqLQq2TrUKCOr0/C1IS2ew/tfE7YIsU357nAvMxug5CiU7c6y5XdQbye9TUy4zFR44HHjUM5FGsb6zZGUmWxYBrf/ntej55NuAvZmEDImxUd5PV0O8n6PBtPjfvSiTPlMS8O5Vva4LOcZCtSs2+fuYrRsmHSSx/AvVT6sGt9VmZGWVeDiRtQ0e442QK/VnRax0LdCZu9/WrugRyfYaXrvW2LhgUfADPYKbR6t8YVPK322SEK5SC2hytSThqFUoNNhBWIZs8LverdRP0ebmE9s3suHJOrzHoez0Pl78eFXMceRyuzdhF9fWUV4H08M2fOSlpNmbdQ5v6Y19Uezoy7xiXfi2fxvT2OJnOlTJZTr4t6jPnxOtyDIJzp+5WxHw5B+l4HwcsKx1HAhJMzL9HrWutwcjHqbzyEOnH82FX3+0OWan2zFWPkeNaPrWe1N+rnytm8er78PuuCx4LOMM5lqau1KXW99HXI14RBda/oZwiFVs5xkyO/bnPZ8httvaLXFbnYnk/WHK/VRtXPP3QDKXJj8rRy+RmHNzQeWt2rjy/MYxInps1Gd6VBqCliuuxmdpbA+fbZMUI63lv6w3978RpI4aVpQx9atnQAeDTBdTGaCGXQEVija9w0wWA0/iAJ6rnO3RoPwlcbkKtemw5iLObl6fRuedC2r6Dr8lRoTsp12cDMog9SbUGX1Od/So5clwTQ5p20qfkAm5rQ5kzB1lp46xdKdHfTnaNkydeXhdg5g/aEpEvTmJiipZqPQfs3Siyo6GSw3IovoYYzv9cxf245kKBcdtU1ocy42vtQCnZCf87KTUXmnOxV4Oezn+MaA+TuLFayvNvTYQwA9NJX+bMHfvXpGY73qVx63LsE+UVe6dp9PktzTBKs7K3xxNY/3s9tE8YYwwQm40JossxPIayKMQauSv4EM+mWNkgK979DWpGfMSEEKaxTNwL5UDupCmNqwaXKOiyfcVkpy19aUWWzNw1jiGP9e478i34QfBcA0cul00WtXU4nMsm1UNNgFZISPAKyB+8ePc+K6+nV7slEwDEAH23RvZMCQWHQeux2F0+SUFeT9u+tT8wGQScdZvAtH5sAGwJXtZYLDfPuciZk8JVqVHy1d0E1LmZzGtX45KmsESwtPSrc6tGrdjWyLzEAYEQIgPM8Jbwwgbvnt+Znu4SeoyJc39AELCtAsDPPGbpwORLl7fi5QF8O3BkgEsNnwU82GIe//jyF8kufxXV92prtamaRyWibrzb8NE5SGxdBr45Q7JJz2iUAyFNpe8f3Ib8OpfrUd4mmSJEHAC08eBtDcdTFjH9SqoP7IU8QwkpGhppA/5QzLD9lVDb6yq07MxPLewW5V4T8qQXPR3ThRjHqYzQTGUyhhGwOcq1qwfEOInOyASHlNjdg3VY24tDf00KmnMfhmRwKTK3E5yJIqXdjxrDwiKlL6ezyupfHVhmaEPUXTgWj6gcfX7E7FMs2PdPdqlit9MlczaPAQLHzUwyWRsa50okBsBNnN/Qxr0QAuDYkYofWzL8c07ZxNDkuzcZlRwliedh/NqR9lgpM3ad3cjUTdGn7HnO+a+d0XKTl0+zN2/js78DafMrYs4/OYvZC2gtKrk1ToEkhIr80X5r4vZQ+NOOZJDc1T3Aexmsso1e7OE1+IWttPbrjp74HJ8LXxVvdHnN7C4c+pfWrUqpF0jt5SvzgB9a4MPJ0uPcmgq4q2jMim8gm+AFOp9nJnoVuDgQY3zVLqXvFte/4Kiucs8cxpbPj35K5BtZycQairNbdni1TMt6wHBMT0+3cLsxyF644dvucGPLqHPrk25eWVtJHYsqzIXJWx68xHlyX/g6XotNkVXpOn8Lw4s89AQ6xxgB0K4tQ1hPaAKYLfjRpOuaNna+eb/eCnS5e7+Da7e5fcTID3ZIu3NRGT88vKUuUipZvZXhqf6+7Tdk1APHFORmSOtaOL0VSn3A1S/PWl/2Zuz0PFKC8wAIyq2kOB9akVhqriG89nqe3GxArqx0gLMH2sBKWpY27FfXsg3HHj9Xw6ecvA8lTUntE02MfpK2qDOb4iJ4bws+UZG+6iygphMzUrR9JNItJ42XIMf7PFKXxTIUNuHQ/XQ9lVZXDvPJ4BzeYDbMA1i530Jp0vG7vE8YztHrYiG//AAAGdUlEQVSsjANgtcYazaw+zl5T4LW30amCSJidd+aObr3PQrEgsZVZN358rudkRVzYIs5ioAFLy6z/V3FsWbg/ylK7mGU7HMG6nyXL3ag1KNyZnZqfrdPyPh6Lu5BjBJo9mTrLcqt5ik1j1HXm3I3qdvRB0AHhjsEXiDoBprpkmkcPjOinG1ljppnsPq7h3foQsopDxwtRygxUHRRyu8UbpKB2vmoRUN2/KssxPUHFWseU15/xN55b2d6sM08XjEp7GAcmEII09HwQiOrTrv0BH4iqQp7QibUD5wE55eS6MC+CGarrvFNmrw7btzEsSdE9+JazIGBhU4NTdUbgFNPCX32vaSBThnXwqeSYDGMh07yG2hW8BwkeA6fkOS81T9O1TD79zmloeqQgv3jTH1hDTCEnmjGF+awodPHsOccZoAEPrQP4Zo2bso/Me+93YEnOia8dOrRC7rA0SD87RitZVKbjMUWYRRi3V1KmHv3pR3mP4CSBwZCacK9jhlygUANIYB1zzgIH1johOOrWYx8Aj+4Pdd2XaH0HBX3y9tOfskMBu+EFNL4+lHvlXfUg3jHpVtXX85kTWy97DwPm4j+dBweh+udZnB3C5HTXKmGd1HdhG6ZkJ8CoKdWqMGQ7PLn11cYOMWNephrR7E677UtF0KsdVpqjAKEbT+gWmUVg8523r0sIQkwtXQIWHa+uUtqbtcNbbAVMhzROW8YIPnE9RqANf0yI2u8p+h7gFk/TwNOYSlYDpZbTsBNCiQIgahjTepe3HuybZ29SCSo8OhL2krfXlgCV74wcEo7QDc0eujeEWl2MLjPB+oZSd8vt23qc9i6gm+O9lKHkVMC97ivuPQJRD9fgUxTyf8Vd1rhe0g312sJ0qzomNUDU6gWjUO4rMMfJ9XF3qtjyskdw2aXi2vAjrvhyj00qIaVLP3ri1YJxHm5M38numH0USg34s0W4xH9L0YpHG8Bp+Cq/Ph2xp+nq00BwAa6k0Creg3/RhwnRTcuhWHYx0d27UGr3nNLItRzKS9mMyBK0CRi/P0IwX7QZoDWX34XUG6Cbzk7SInWqo/ejTay0lBG13kEaEcDTHcB16fL6geTM3F56CUSeQrOlpR97YZ5HDjzm7mBHqQPIpu8r56eYAh1lXDhqsoBcexNdlEhoWWO69W3wc0BBCtsK4McTsxH/+Fsaj+WtS1962qN0DwqHWd0E11yeiO9S8MweU4PlMTT9sB8ir379DineSopAQ8q0eXdXtJZf0dmdjfZHk5l5iWMeL4e3clav5KM2hDvuvN/7//72c+lf93vi5zo7w7vxgTgTR86O+d07SinOe+r8pY4Ha9BPu7Rl+Q4wj/wmk9B/ZyPnbcwE0h792QIo+TYpMxlXMMPQ6bqTch7HAtS/7uNv6MhLc/ZHKdc7/96pMEUe88YcGsFuwR6EgtHTGg9PJxq7IX4JDV2+5mtbcVZ7UUOmo9nNGIpJ+6ZfH0/PLvXRrRsFpMrwRNTLoBch6KlJ0PQTaZUW+aEi2ZUHAM5TfKpJ3eEoIztQwqPXBZITbv7gLU8boNCUatcrNcphUVY4oB7bKDcjAVTHOxmmL78lh0OWyfF4efbxno+cdo0pfMpXTJvKsImacPnA5IwHISm3TwqcRCubRBm9OWoi2vs68RJwpT4uQl96HfK7grAGDOtu/SFkue9L/7P//tf493/5j//84/7nv3ytf/q3Y5Fs1zM/QbGngFSZv9AKPm3QzDzLrR1uuZcOV+KOnxykf0ePxlFs9Y/8SrvY4YnJVMaKK598xaXbKE4oc0dqR2bmiitTT4TqNyW7y59P5xoUJT1T/FToXXkHr8CNCy2+570EMEgp7VjxlbiHThPH0p2TIny0vMcqKnqfRcl+dhvlyNoXgt1ZFvWLtJ922F3MbtGuO6ivlcQcaenKWmrYXOVMS4qllT5WMBRLV3zlzncQaElbq9ag98cciQ57gfnoHUtXLl015rhSWWIGC5Sj/a74Ss+zTnTda5L2AOPSV+5m0BJIWsS0k3qQrScys07S60LF67fvZYz8ku2o13buPnsI+U1t780lv4/eUa0G7iQPVjJ29jFpXCBCoUdv3fGdbmodVlSvc2jnO2puwf4e8+eerPuU/G49gXFb8ZU2en6t3EvMR8tv3d8m6jJi15hIy29UPrLlV9awrXcs3XvFHdX8+gl7XPnOP//6v7/++7/+H6vpvl06Wf67AAAAAElFTkSuQmCC"}]}
