{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"#ffffff", "background-pattern":"" , "items": [ {"x": -783,"y": -168,"w": 3111,"h": 1837,"type":"image", "image":"jpg", "image-data":"/9j/4AAQSkZJRgABAQEASABIAAD/4gxYSUNDX1BST0ZJTEUAAQEAAAxITGlubwIQAABtbnRyUkdCIFhZWiAHzgACAAkABgAxAABhY3NwTVNGVAAAAABJRUMgc1JHQgAAAAAAAAAAAAAAAAAA9tYAAQAAAADTLUhQICAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABFjcHJ0AAABUAAAADNkZXNjAAABhAAAAGx3dHB0AAAB8AAAABRia3B0AAACBAAAABRyWFlaAAACGAAAABRnWFlaAAACLAAAABRiWFlaAAACQAAAABRkbW5kAAACVAAAAHBkbWRkAAACxAAAAIh2dWVkAAADTAAAAIZ2aWV3AAAD1AAAACRsdW1pAAAD+AAAABRtZWFzAAAEDAAAACR0ZWNoAAAEMAAAAAxyVFJDAAAEPAAACAxnVFJDAAAEPAAACAxiVFJDAAAEPAAACAx0ZXh0AAAAAENvcHlyaWdodCAoYykgMTk5OCBIZXdsZXR0LVBhY2thcmQgQ29tcGFueQAAZGVzYwAAAAAAAAASc1JHQiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAABJzUkdCIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAWFlaIAAAAAAAAPNRAAEAAAABFsxYWVogAAAAAAAAAAAAAAAAAAAAAFhZWiAAAAAAAABvogAAOPUAAAOQWFlaIAAAAAAAAGKZAAC3hQAAGNpYWVogAAAAAAAAJKAAAA+EAAC2z2Rlc2MAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABkZXNjAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAAAAAAAAAAAAAAAAZGVzYwAAAAAAAAAsUmVmZXJlbmNlIFZpZXdpbmcgQ29uZGl0aW9uIGluIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAALFJlZmVyZW5jZSBWaWV3aW5nIENvbmRpdGlvbiBpbiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAHZpZXcAAAAAABOk/gAUXy4AEM8UAAPtzAAEEwsAA1yeAAAAAVhZWiAAAAAAAEwJVgBQAAAAVx/nbWVhcwAAAAAAAAABAAAAAAAAAAAAAAAAAAAAAAAAAo8AAAACc2lnIAAAAABDUlQgY3VydgAAAAAAAAQAAAAABQAKAA8AFAAZAB4AIwAoAC0AMgA3ADsAQABFAEoATwBUAFkAXgBjAGgAbQByAHcAfACBAIYAiwCQAJUAmgCfAKQAqQCuALIAtwC8AMEAxgDLANAA1QDbAOAA5QDrAPAA9gD7AQEBBwENARMBGQEfASUBKwEyATgBPgFFAUwBUgFZAWABZwFuAXUBfAGDAYsBkgGaAaEBqQGxAbkBwQHJAdEB2QHhAekB8gH6AgMCDAIUAh0CJgIvAjgCQQJLAlQCXQJnAnECegKEAo4CmAKiAqwCtgLBAssC1QLgAusC9QMAAwsDFgMhAy0DOANDA08DWgNmA3IDfgOKA5YDogOuA7oDxwPTA+AD7AP5BAYEEwQgBC0EOwRIBFUEYwRxBH4EjASaBKgEtgTEBNME4QTwBP4FDQUcBSsFOgVJBVgFZwV3BYYFlgWmBbUFxQXVBeUF9gYGBhYGJwY3BkgGWQZqBnsGjAadBq8GwAbRBuMG9QcHBxkHKwc9B08HYQd0B4YHmQesB78H0gflB/gICwgfCDIIRghaCG4IggiWCKoIvgjSCOcI+wkQCSUJOglPCWQJeQmPCaQJugnPCeUJ+woRCicKPQpUCmoKgQqYCq4KxQrcCvMLCwsiCzkLUQtpC4ALmAuwC8gL4Qv5DBIMKgxDDFwMdQyODKcMwAzZDPMNDQ0mDUANWg10DY4NqQ3DDd4N+A4TDi4OSQ5kDn8Omw62DtIO7g8JDyUPQQ9eD3oPlg+zD88P7BAJECYQQxBhEH4QmxC5ENcQ9RETETERTxFtEYwRqhHJEegSBxImEkUSZBKEEqMSwxLjEwMTIxNDE2MTgxOkE8UT5RQGFCcUSRRqFIsUrRTOFPAVEhU0FVYVeBWbFb0V4BYDFiYWSRZsFo8WshbWFvoXHRdBF2UXiReuF9IX9xgbGEAYZRiKGK8Y1Rj6GSAZRRlrGZEZtxndGgQaKhpRGncanhrFGuwbFBs7G2MbihuyG9ocAhwqHFIcexyjHMwc9R0eHUcdcB2ZHcMd7B4WHkAeah6UHr4e6R8THz4faR+UH78f6iAVIEEgbCCYIMQg8CEcIUghdSGhIc4h+yInIlUigiKvIt0jCiM4I2YjlCPCI/AkHyRNJHwkqyTaJQklOCVoJZclxyX3JicmVyaHJrcm6CcYJ0kneierJ9woDSg/KHEooijUKQYpOClrKZ0p0CoCKjUqaCqbKs8rAis2K2krnSvRLAUsOSxuLKIs1y0MLUEtdi2rLeEuFi5MLoIuty7uLyQvWi+RL8cv/jA1MGwwpDDbMRIxSjGCMbox8jIqMmMymzLUMw0zRjN/M7gz8TQrNGU0njTYNRM1TTWHNcI1/TY3NnI2rjbpNyQ3YDecN9c4FDhQOIw4yDkFOUI5fzm8Ofk6Njp0OrI67zstO2s7qjvoPCc8ZTykPOM9Ij1hPaE94D4gPmA+oD7gPyE/YT+iP+JAI0BkQKZA50EpQWpBrEHuQjBCckK1QvdDOkN9Q8BEA0RHRIpEzkUSRVVFmkXeRiJGZ0arRvBHNUd7R8BIBUhLSJFI10kdSWNJqUnwSjdKfUrESwxLU0uaS+JMKkxyTLpNAk1KTZNN3E4lTm5Ot08AT0lPk0/dUCdQcVC7UQZRUFGbUeZSMVJ8UsdTE1NfU6pT9lRCVI9U21UoVXVVwlYPVlxWqVb3V0RXklfgWC9YfVjLWRpZaVm4WgdaVlqmWvVbRVuVW+VcNVyGXNZdJ114XcleGl5sXr1fD19hX7NgBWBXYKpg/GFPYaJh9WJJYpxi8GNDY5dj62RAZJRk6WU9ZZJl52Y9ZpJm6Gc9Z5Nn6Wg/aJZo7GlDaZpp8WpIap9q92tPa6dr/2xXbK9tCG1gbbluEm5rbsRvHm94b9FwK3CGcOBxOnGVcfByS3KmcwFzXXO4dBR0cHTMdSh1hXXhdj52m3b4d1Z3s3gReG54zHkqeYl553pGeqV7BHtje8J8IXyBfOF9QX2hfgF+Yn7CfyN/hH/lgEeAqIEKgWuBzYIwgpKC9INXg7qEHYSAhOOFR4Wrhg6GcobXhzuHn4gEiGmIzokziZmJ/opkisqLMIuWi/yMY4zKjTGNmI3/jmaOzo82j56QBpBukNaRP5GokhGSepLjk02TtpQglIqU9JVflcmWNJaflwqXdZfgmEyYuJkkmZCZ/JpomtWbQpuvnByciZz3nWSd0p5Anq6fHZ+Ln/qgaaDYoUehtqImopajBqN2o+akVqTHpTilqaYapoum/adup+CoUqjEqTepqaocqo+rAqt1q+msXKzQrUStuK4trqGvFq+LsACwdbDqsWCx1rJLssKzOLOutCW0nLUTtYq2AbZ5tvC3aLfguFm40blKucK6O7q1uy67p7whvJu9Fb2Pvgq+hL7/v3q/9cBwwOzBZ8Hjwl/C28NYw9TEUcTOxUvFyMZGxsPHQce/yD3IvMk6ybnKOMq3yzbLtsw1zLXNNc21zjbOts83z7jQOdC60TzRvtI/0sHTRNPG1EnUy9VO1dHWVdbY11zX4Nhk2OjZbNnx2nba+9uA3AXcit0Q3ZbeHN6i3ynfr+A24L3hROHM4lPi2+Nj4+vkc+T85YTmDeaW5x/nqegy6LzpRunQ6lvq5etw6/vshu0R7ZzuKO6070DvzPBY8OXxcvH/8ozzGfOn9DT0wvVQ9d72bfb794r4Gfio+Tj5x/pX+uf7d/wH/Jj9Kf26/kv+3P9t////2wBDAAMCAgMCAgMDAwMEAwMEBQgFBQQEBQoHBwYIDAoMDAsKCwsNDhIQDQ4RDgsLEBYQERMUFRUVDA8XGBYUGBIUFRT/2wBDAQMEBAUEBQkFBQkUDQsNFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBT/wgARCALRBQEDAREAAhEBAxEB/8QAHAAAAgIDAQEAAAAAAAAAAAAAAAEFBgIDBAcI/8QAGQEBAQEBAQEAAAAAAAAAAAAAAAECAwQF/9oADAMBAAIQAxAAAAH6B9vg06yUkRjQiCxAIEFDJSFZjYCFQiAQUIgAAEgFIAASAAAqZiCIYCFQCIFBiBAAEFEFIYhwrAAVIAABQIVgOBWAhwUhwAAAA6JQYCGADlYDCGoJGAKDCAYACsAAAAYKQwUQVhDolYDlY4ag4asylF3Z1quNO8pMQpWJEKkgAgAY5SsGQBUCQpICoAQAIEAEFAgASAxCpIAoCArAQAAAFIBIDEAAACoQhUAAAqQFYDlBiAACiGogADVwgABgoMYZNRQYAgNUMBwDURDVgACAYDlBiGAwlag4YKxjlY5WrjKGu6beZo3lUSKlYkBCCxAADgVCuQVAgECIKAFYAIQwEgogKgAAQkACgQCQBAQAAUgFYAIYhiABAgoFEhaBIqQDAYhDAAUGIAMoYlYgGADhyg1AAAGAAMIFaAArAcKgAHKDAAAY5SVgMFDKGrHK1Y4cu+beZp3lCRUkVCAhBQgASsRjYICCgQAIYhWCKgFEBAJGoIEAFQAgQAQCsBAAAgIVACsAABAAAgqGJBWJFSGOAKQwURArAAhgCsYgABjlcoAwABDABhANQYAOAAUQogVgAAMFcrgAaiOVjVw1ascEu+byzNOsqhMQpWCIBAILCGooY3IIAEAUkFEQAKiQoFYKIBBakAAQAiGIKBIgClBYCAEQAKgBWAAAAIAAAEgKnDVAADFRAMAAAVjCCgQ4auUGAStFQogoA4ARqDURyiCgAgAKwAYSg1IYxKxhGSgxysFcOXfN5ZmnWSkiFSCwEgIBDAauMLChEIYgABCsAAQAKiAEAChEFAgASMQCoEgIAEFiEgMQh0hDpIAAAAgAAEMAAAAAABgoADCCDVAkcrUGAK4VNEoA5BQYAMFIYxAgCgwAYhq4AUHAMBq4ag4YK1yDN3Z3nGrWMaEQBZiFogmIAZSoyXPOtO8CIKDFGAKkAEFAkAAQxAAIgsIKVAQqARCoEgIQAFAkSAAKiCgVAAgAAAAISNQAAAAYACgwgGAAIcrVgA4FAAAABgAAOVgAxAMAAYAErBXAAwAauBWA4DJoGEdGN5S6tYQUkQCCkFiQHKK4zmspdHTkgEFEABSAEBCCkCAAAAAgQMbCgIKBCEjpCQEAqBIIgAAUQVWFAgAAQUABIhjAQAMJSnIrWEAQU4YAoCsBwKAAAADAAGAK4YAAgAYDAJXYZrUABgCscA1AGEZK1AN/PeyXTrAY0AJEAUAiHK1yXPOg0dOSAQIAAgAKQkAAQACFAgEAIkKBAFIQIlLABCQFQJECAAoABYgoAAAQxCQBWCAKxBBTgAYQAA1AGoAwgVgACAYAMFARysAAAABgoECuGAxDBRHKDAag4YK1BjN3PpsjTrCABUCRDAQDBXGU1kad4QUkSCgDEgIApICAABFRKIUgECIEKVAhIKBYgEAgsQgEgADBUAUmSiVqIrCAVAgGADgolEAgohgogoMaiCuABqAAAADAFYQAMAUQABqIK5QAHAAwUQGpDAagDCGrVgBvxvZm6dYBAKgSADEAjJXLlKjXrCopAgAAoiBAQAKwAQAAIgpAIBIUgsQCAKBAiAVJAAEADEAAIEFACkCCKkMYBBaBDgEMAAYDUEOGA1AAYAAAoMACGCiDQMESNWKGoAQwAAGAK4AGMFYDlagDA3c97ZdOsiIAoEAhgIEa5TWUY2a7kpAAqcFgAgBEAAIKSACABBYgEgoKxBSQAVACgoRCAAsSgAgogAgAAEAUkxsY5QBgoEFCAArhDGAAA4agAMAAABXAAwAFAHBaQI1ACABgADAakAAMBqAMJWA1Bm/G9mbp1gAQBRBSAcKg2Z05dmdat41awlEAoAQAAWAgQAQgsQAAhAKwAQAILFQiEAAAWIQAIACiAEBKWMUpYAIQWY2NSVgABAMQwAAAYDgAFYDAAAIYKxDAFYkaoY5QcKiGIYAA1AGIcMBDAYKAMJWNQBm/GtmdatZBIgAACiABrlLnNZZuNmjpzQIAAqAgAKVCIEBAIApIAIBCoECACCilIUkYgEFJAQAACGAgAACiFSQCsUY5QBAMAAAABqDRDgGoAwAcCgIKDAABWAKQxwgGAACiA1BwUQwAQwGAKAMIag1Bm7Gt2Nad5BICABqAIBmedBtzpHP05LRQAAIANUiFQgFIARAAgpAJAQUCAARAAqLEAkQCCwEADEAxAAgGIVCAqUMBiAAABqAADAACAYAAwHAoMQDABgorgCGAAoAACCiNWEAxAMAABgJWMBysFAOjGtuNatZVAgGAhiEMFylZnmi6tYx1lAAAIYCQEAgpWACABAipiABICAKQkAAVAkVgIBWAACiAACiIAAAEKxAMAAABRAFBwAAAAwGoADFDAAGADAJWoOAABQAGIYDEOAYgGAxAAxDUQVgrgVjA341uxrVrKFQAAACABhKzdjezOtO8aN8wAAKAEAkBAKikgCiAgRDEACoQEAhUCQABUIqEQhUAMQDCAVAIhiGIQrAAGEogpRAAAAwAFEAUQVgMIYAAxDCVygwAABWAAADAAhgrEAI1BIDAFAAYBKxqwN+N7cXVqCAKIAAqAABy7M6zlymtWsad4SAxAAAAqQIgpBQACBASCiIYCCkAkBBSECAgpCsEQAADAAEFIBiAQJjYSsYAAAA1EQACsQI1EFAAYQAMAGrhUQ5WMBDAFYAAhhDUAYAAAAkBqAMAABwAuSgHRjWzG9espGJWIAQUQVDQXPNymtk1hc8/TmAgogoCIBUCASFACAKQDEJAARBQIEQCoEAkQUCsEQAAAAKICGIVAxCRAMYhgCgAAACAKxAADCABiGCgwHApAMBgoMAAAAIBqDAAAAAAQUAYDhAA1FYwjfne7GtWoAACQAAAAHLlGS55015enIsAAAEIEKBCAAEhSAKAECACQEFAgEioEJABUCoQEAxAAAACRiFQMQkagDAAgAKBAEMVMAgAAAFYIDUBSGEMBgoA4AGAACgAMAABiAAGIYhhDAABWrHBLuzvfm6tQAQxAIYCGJMlcZ51kqNG+YgAgpAACCwVCQABAhSAAFQAkBIAKgBIqQCBEFIKARACCgDURAiAACkJGrCCgIAAAAKIAGCiAAoCCiiA1IYQDABgoOAYAA1AEMBgAAAgAAABhDEMFBgrHBLvzrdjWrUKIKAEAAAAMcZ51uzvGzn3zxsaJREFogqQABUkAEAAJAApBQIARAiCkArEIAEgFKlDEFCCuCwlBWIARDEFA4AUAYgQAQAMFYgGiUABgCgBDCUBGNUMYQGSpGoADBUjAJQABCgQAMAHAAAAK1cMIF3530Y1qsVAQUIqACAKAHGUu3O3Lz9OeFyAACogChAQCCwEACAQICCgKBAiAVgIQIqBUQkAFQAAA4BUAILAQIKkBq1QIwUEyAogCg1BDRKIDUCAKBwAOCiUAYDHArAYAEFADlAFRDAVCAApAjUAYCGNQcEoBuzvpxvXcoAABUAOEKx0QUZuya2ZurWdW8ggABI1EBBYgABAioEACQAKQCoAQIrAQgBEKkgoCAAogAAACpWADUhWA5UFCOUEKwAaoYAACGAIBKwoCCGAArABgOBWMACGAKAAAACGKxyoBgA1EaggGEMIagG6b6Oe9dyhgAgAAASFEFEZNZ5rNW842IBDAQDEiChEACALEACAAEhSpwqQIhIUgECAqAEADAAgpAgIQBTgMdHBDohUDgpAAUQgogCgEFAHAAwgBQYAAwCGrURgEMFaJQABBQAAAAagAMACCgIYQ1Bgbpvfz3ruQAAAAAABAAILlLnLhZhrKoAAEAAIARWAAIBBYQqAEAAJClSBEioAQAIEAAQwABqhIqBAgACohjVAgogACpwqYgCkOEMAAIYArABgAQ1BgNQJGoAK0ABQAEMQAgrAAAcNSCwEENWAwA3TfRz3quQAVogAcAUgEAAbJrPOsbMNZxRUIKkKBAAAJEOxAIAAQCsAAQCQpUCRAgIBUAAkagwEAAYoBSAAAxTJQAABDABICGFEFIYQKDEAwAYQwAAVgOUQaYIArAAQUAAABAjUGEAwlAGAkAGoAwHLuzvfjWvWRQAkLRCUBCkACADJdmNZyhq3nXcoACkhQIAAQrCQoAQAAgQVWAgEhSCkgAgRAKmAhgAAAgEKwgCgBDgCgQAAAIAQUAAQVgAAMBwAogADUGpI1ABQBgAwEgrEMQAMIBhKAMAAYgABgA1cbpvfz3ruQVEMAAAEhSAAEM243nNZRp3jDUxQABALUBAACRAgrEFgIAEAWIBCBClQAgEgAAAAAAoKxICAAAQWEAUQUBAACpiABgIYAAAOUAAAYAMJWAAoAwAAGAhhBRAAxDhqAAAADAQDAAGErNud9ON67lAMQxAACCwEAANduNuMlxsDTvGKMQBSASFIAEAxACCJSwEAkBUCASFIYgoEIYAAAACBEKhABDEJGoNUgAAJGAgCgIBgogCgDAAAAGADlFYAgoAwAcAqAhgKGFEojUGIYAIYBaIQDVwgGBtzvqx013KQGIAAAEIKAAQ42TWUuUuUucujeNG+YACABUrAAEAAAkAFQgIQIgoAQgAKEVIBgIBgIYhJq1nRrGjeNOsaN41azlLuzrbne3Ot2d9GN5SgwURI1xQABiGAKDAAGACABqQxGSgCGAAMcCkFJGEAAAwUGAUBApYQ7VDAIYAADA3Tp08t6rkAAsAEAAIAEADBdkpGc1nnTOfpz16ygQAQCoCxAAgAAASAgsQCABWAqIAFQIBiCxGu50bxzb56dY1azzbxr1nKXOMLENc416mKZStcUzXdje7Otk10Y3uzvdnThDAAVgADAFIEFLECuGNUMBiGIYDglEFAChCGIYWuEMACiGpCpwBRDAAGAAC7s76ee9dgACQBC0RKAgAgAAMlQ5dmbnNI5unIoEgoiABBYAqsBAAAAgRUIgEAqAASFI06xyb56t45989Ws82+eFjEMFSZzWu5a7prRrBG6a59YyVxq1NkIxGBkYJku7O9mddOOm3OujG+nHTOUBWgENRAGhENQYwABDAcASgUwgogAAAYAMQwBSCiABgAANQBhBRLtmurnvXYxCASAWAKhiBAAAAAF3Y3szpWc3TmkBBQJBREIYAY2ABQAgAQIqBCQNG8cu+fN058u+WneOfeMLnJQBDEAGUuFm2a0az051zaz0Z1osZtl57nevNcb5rRc7FwTJUA0FQ0RkuKBszrbnXTjr043uzvpx0343kqAARqDHCGAgohysQDAAGIAGABDUABgAhgAArAAGEoMQG3OurG8LAQCAQBYKBBQgCiAIlBm7G886xs07xhcgAFIBIAAgEFEFAkKBCTn3jj6c9G+fPvnx9OWjfPCzIxTOaVMxQGuJka7NsumzdNarnfnfPrG/OtOpuzdNm1cUYGnWdudc+sbZdNm6XRrO/OtOs7s612ZS42AzGsoxM1wTJQxsyl6MdOrHTPN6ufXrx06sbzmiGpAAAAwGIAGAKIqcAwlYAAAAAADUAFaEFpAMAA2Z118969QABCAAEAwABDEFgCEuyayzc5dG84awCAAAVAkAEAAY1z758XTlz7xz758fXlzb543OS5xrsyMQMlSChjZlGFZAYJumuXWOvO+XWd2arcE6c64d8+3PTj1jtzvCzQnRLwb592d8OsdMumzE3S8msdud8us7s6VYpmazNUgCgI1RnKrCMlwszlxTfnfTjptxvr59OjHTsx03Z24BhRDUBEA1QBY4JWMBAMBAADGoCuEMQAMBgbsXox1wsSFAgEAAAAAAACCiQM5rZnW/G9G8c/TmACAgAQVjZzbxw9OPJ056N8+Xpz5N8immyaSYWZLhYAIzhqgMjXc5zWFmKbpeXWd80k02ded8Wsb5rbLwa5yOevLc5G+Xh1juztHFrPbmxvTn342LGb5d+d8esbZdzXBrn3Z3pswOrOuXWdsrNdm2a12BnGNZSiChkIDKMayhqkyNdZ5vVjp0Y6bsb7OfTqx16ufTOUABiABgNRAAAAEMAVgpDAAAAAYG7Ounl012AWJRFQAAIAABgIAADKOnn1251p3jm6YxsEExNG8cPTlxdeXLvlx9eXNvmq2mU0JgZGNgNcWVQIDOXKNdhWUuqzZCrTc75rVZquerOuXWXHTN8OsdM1vli985LHRrGb5SWOokfvnI46pI/WJDO+XWcU6874Nc862yxu8d2dZrG6xIZ2k4tZ7s7wTnuezO9VarnpmtNiOjOtdiTZLjQMcKnDARnLjYGyXEVEYmzOu3n16MdOnn06sdO7n03Z21YAMQxDhUwAAVwDAAAFILCVgbc3p59MLEABSGIAsQDEAAACAZnnW/G8o594hPT5eDvw498uXpzx1nTrGxcjWMZiFhGFioAxsUMVBtzrGzFM5VWq52ys5tZ3S5y8W8dGdbZY/fPqzravBrHTN9GdcGsbl6c3l1BOmawTi1mRxtEfvMhnSIrfOVx0aQu+cnNpInWJXOwjdZ7prZLH6xvl6pri1lx2zXJc4V2ZuqsE3zWJhZsjKXGwlyTGgylYCTJWIcrADJSTXWqs8unHTu59enHXp59O3n168bylAAAolYAMAhqUQBBQMI2y9PPprsAEMQAAUgCwUQABHPvnH9OXD148+8aN8+Hryxud80rAcY0kahjYgBMLBWmBjZkuRgmcu/O9Gs42bs6ws0XO6XYcWs5nTnXJrOu57cbwqO3zkcdMiN1jqmuiXTZxXMlnYRG8S+OjI3XPvm85RIzWJPO0RO8SuNhyazo1nrmsEidZmM7CN1jqmt68zPOSU1gnBZ1y9C8VyHbnWqtNm6XZGiwOmXVZibJWYIG2XGiXIyAQ1YQjIyhVibJVWhMl6cb6efTpx06efTt59evHTdnTVgA5WEKgYQAAG3N6MdMLAAABDABBWNnPvEd05cnTlp3jn3y4uvLG5yM1cKkAjGxAhShUI112IaJddyzZNabnJd01lHPrIdGbo1NVztl3TXHrGNnZjeFnDrn0ze+Xns5NYksdBIzeeiXqzpVDaxN42Ly3OiyQzpkRvEvjYBEb5yudix9xuXqmhILWJVVWlOAlVCNudsvYuBG3MhnW5eS45yRmmvHch351qs02ZR1zXLZim02zWqxG6VCQXbLiiUN0qpQGQkFKcZKhGyG0kahy2Yx1Y69fPp28+ndy69/Pr0421cADUEgom2Xp59NdgAAIVnLvEf148XTnydOfF048vXkjtzrdnWzO9es69YxQoMbEYo1SZGFIEyjToJlKVouVZumsEwTa1053rs03ORvzvRrGi53zW2a5bjRrPZneRxaxrskMbDg1kTum8UjdY6JrrmkkLrMtnW1RIPWJvO0MhtYms7IVQ28TONhjUJrE3nYmgh94lZSuJNMsjWUR9mKyIRHWZEhKqjWdiyEuJw3OcvfNYHLrLjtmtSaNQjsmtSa6I65rWY2KN66xAbpcBgbFxGEZKDGIyVyC4oUGBpTZNb8dOjn16cdOzn0kefXu59Nk05Bdmb0Y3q1nl3iN68Y7rx5uvLm3z0bxp3nZJums5REOss6a5S4XOvWQRjcisF13KM4DRrIZy5nNrKNkuZy6znL0Z3ul5tZ12bpdsvNrPPcdE3ul1WcWsdU1vmsEi98+zOumaRFa59U11yqou43NdsC8NmtJKVrqSJ1mazpDIbWZrOhQhdYms7cKoDWJ7OgCD1O6zYER1ZEgYxxWaCUVGhOGWVMjVXCz3TW81nFZtjumknDYzumsjiuWbl3S81ijNeqXQYWZR0zWBhTjMyXWmSs2S4I1SZqQKxIwUGA4DGsaxjCa351046dGOnfy6xXfzcHXjlZ0SsYwHKqSBlKrEBnNbJcDVrmLsl1aziiNk1jZquVZnLnLz6zhYzfLpsxNkvVnok5NYDpm8o5dZ59Y6ZrdnWNkbvG2O3O1XFcaLJLPRpgQuucrNbmkkXc5ndKGFkKT7RDIC4nZrKVmqyKsmZoHLBb5zeNliIvWd8vbKW4pXLmaoRERHZXbKrOYjyYBRImOyusZxmlJXO8jWcVmadjTTisSdedb10JpsDszpVz2ZSs3y6LMRnTnTXTYka9ObqpIVnm7FwFYRtlxrFBSM1Q0VuUoCIVOXu5dt0nNvGNjMoxBVY4KxAE2NYIhm/PTZm8HXigTdNadTWyjYbJeXWcLA6Jca57nZL056bpdNzzXJXXnYc2saLnozrdNKo3XNJIzo412ResdS9WdByXMdczU2zEitZ2xIKhWV5LDNZAYJBk+oKIPWZReiVqJX7iwTaEiqBSfmmKotnmuZCnKVAxMpstE1ywsTtjpxxHOSoKEYbCSla6E47N52Shy2aU6ZrrlVcVyjqzroXWnPYk6ZvZHPZrscdc3lLzXKojrzrJdFyVlL0Z1imvUSOXfNYJhY1I3LgFAS5r2cum6OLpyRjZsmma7ECbJca1jFZvzrXSMo2zWNzzaxrsVbZdkc2s6xJ0TTOfWSXdL2Z2jk1jVc7F6c6Rx6xqs65vdNJODWOayRm85RI7WNBKzQKou4RJTTMaiWdyyACIRO87FAK+k4bLSAr1zYppqIFeubBNNQxSus2JpgY1VmZ3WWMwK/nU9rOYGqISanrnKspdRExLm2ka4j1kDqlVmg4bOuXqhroTls3S9qtedNFm2XumnHPZosDuzrJea51oL151tXmswuSXol3zXPc4hW3N6JdFmIGUvRLq0xAcbmsDs59d2c8vTnqpiTZNM03Iqs2S5S8+soLN2dZy6bMpdO8ZxsXTZz3KTfNbDA5tZzl7M72Shw754WdOdbZUcO8arOvOt0ovJrPBcd010zSNVzE6z3y9U0KrIO46ztVARKbSRUA4E4yaphLhZXYslNSElbSx2gKJW0srTgpJCRIV1qCONIe5mazhVqkgs2f3M4K1kDjU3rOymIic3dUkguRwy86zhlAca8bPWvWM0JxVmSM1lGJxXIvZLulK4UVmyOybDnTVch251ta0M6LA3TXZnWBo1AZ1Z1nLzayAucdE1prCzt5dWzo3jbNaLnFMazjom9bOjUSFb86DmuVQdGdb875tc+TeUm5d2aq5bkN8115201WcNwWd2ejER2+eq57c73SqtNkXcdK9+dCoitY1EvNCC6rIK5mV2iBIg2ElaQGuyty2azIFRXZJmugYKkrEWigBrV2bMrAxrFK7FktAElZymd52CMLOaWOzqd1jJQxILOpSzqsSZLwyx+bPamwFwSMmuqO+zEZHrzEgnQNcY4KEkprIZzGlNy9sucuBx3Ks6JeqaI5bNVjTszvYutOewMjszoNNawNkvVNI0UhJ28+3RnPJ05tejG8jRc69Rmcu2VJx7zruRemayMTkuQyOmVGizm1jdNd+OmconHvHNc7I7JtqkjdY0ax353tlDGojXPIk87ArQQesSi9UoBxJGXM60wFULmbNSTViFZVsasm87BqzBKvm2jUasDlSJiwGNogVtLGuQlSBWZLNa1EDWlWiw7yxQVG5urOpjpglBkJnXdZ3WJA1rB43L2d9mKhzEfmytm8KxI+NEspW8YRGqiRjdaRqs4kJZA2LnLy3PNckvfNbZXXFc4q47prbKk5NTGA65ra1inLYlZ0S7Ze7l225nJ05c2s4gvRNZwjl3jFBeiayTE4d4xTZNdmd5RhZwdObl6M3tzsMa4N89Vz1Z30zSEkZvnqSQzvcqEkZrGiyWzvNQxSH1nRZNSgUoiLMUl1QVikRDqWBWIhI3VKAjUICTvrupysRXUmq6VIAK7cza75QSFV+WXTpC0EkBHRc9eojAzIbGt9S1gMIiJpkrrLhgRGdJZuxmNKI1dMTVmSkKoyNSy5sMgI40x3L1oKJH2azolkJrKMbI+51GyakZc5ROLU1jl75rdKHLZosS9WddKs5rNVnby6dOdcvTl0505cbOPeFBZ0TTgrj1nWCdmd5AaLOe5dSGOmcKsUjd80vdNbJUiqK3y1khNbpREcGs8JIr0ChVoSCslDrCkCQEdiyNgIVQ8jWXsQAnIsJjdm6YBCElUxq17jGCiVPK1aZANQgo77O5WJAwKpjVr3BRkMCoY1aenLCwUAgOe5nU7DIAIzOuQm94AHHJNROdWOzdQONaw0uVkwZgmJFTQTk1sMoa8UcGp0JICQNJxG+WVzvarMZIzU13OZI51kBxWazdNSWN7ppxzanHrOFZHbm9vLt2Y1x9OfHrGNiTomhBea559Zymu7O9soYWR++YdmN9Od42Byaxw7xtiSx1KSIiN8tWsyeOmwSI57IfWe+WRmiMbFURcc2pMS5GJjZrK7E/W8aqMdSHjBJewGI12VHn0uXTIgC4pCRuqUpGUNdVzUsat2jMTIRCyMl7Q1pkBT+erZ0zmqMUaxURMkx0xmKXEyqs8uln1NyNcBnDLGZsrW7WWJXcwWOk2dKbrBdGbyVEZ1N2NNtBpzrl1OrN2y7TopEXHNcyS6M3os6KxWGjuJaajJZBM14iG1iQmu+IfNm9ZztiaxmZvHTY1EJOhbFaxtxru49av14TOd7bK9vnqxuznBrMZrnP47Kyr6x1Y3YLYbXPmiem8Co3EznpNXMPrBnU21x3NOksqyOpD6xz53P2caUbGrlp0Jw6yY3ObzGpROe79vOVkHHTNTW8Rp55w7eh9effrNVxqSqU3iHzaHw7+l9+W+5p3PpYN579Ygc6ovm9Pqfq8u+qTx6W7rjo1K1z1VOHf1L1eZ155w6+g9+QU7luIxv0jvzzSk8ul168sCj8euk9D7cwonLpfevMPP8Aj0zL725Fed+ft6P34o8x83ok+nK/dsYR595+3o/o4o8s8vonevG9dc80tH49PRO/FL5T5u8905X3pI/Nq+NXfpzwt8u4dJvWfQtyNmq/Ja9TNfPcJOy8Ww81CyWinbRszrsvLUPLw3M7LjbR5ndF6a0LzWdK7pavrmi053rXWm4ctYuMLLDnpIzSMjSkDrONklndl49uzl3hunKM3ySzedqzBNi8OsQO+YtlxvRZquemawSp75bJq3Y6cus6NZ65WtIvPYXSb5LIlmRqQlolzyJfWkVy5mFkKomZBx6dtvKZlMakpqV3Kg8t+sdsdpSs6kbJfeYvLybh29j9HKRsqvPWFtj6Yj5PGfL6PXPTysVkdFXzbf0zxHlXm7Xjvzt+sso+LetzgPOudkbbzvPWlUstc1xFJiPY9Eu+sqNzbZeWq/nXn3G+td51EBlIkhqQ6+P+Tt7B6uHdqR2dRPPVx68+BfJ/N2vXTFj640S1Pj0vvblzV5vx6TCWjc6tSo8t2zWd+lHxrnZtizG1XzemJ7UgiDksud91RZzSWS64tZqExd2o/l27OnOPJHOtupRmbNc4cu8nrGjTHGpTUrWueSWXHWtY3OdOeEu+ait84nXO9461Pl2k9Ykq0TerfPRjVp59K914dM1njpssr9zx2XeyA3z6JYvO5HOsbmlpctM9Y2EcdPPt23NCzcbLt15aqxSPx0lY0HmfPXpPflvsdVrGpHG7DvHm3PeFzfu3MqPiK59LXqQyeV+bt6j6/NK6mop/LpZrZPefK/L35rn1f1efRZD5vHy7Wztzj5PEPne72T6Himd51FD4dr71xvs8y8nePs9k9Xn5batz1I6zNabk+fPF6fbPZ55euSWtXNrmuso+LTsvbOs5CtJ3E1c5nhHl7+idF068uFaJzt77c+tKjy6eY+P1++e/x4y0bl0sHbhM6mJ4x4vZY09Q9PGMlonPXoXp8+whs78g+f7vYvV5bDuVPG+nrxm9QPO+Hbh49fXe/Himq5rFi6c+hYyPNfL6bUeh9JW009eE7TKdz6QPHt6BUisFvl2dOUssaee8Oy59PRdOzU0dePTc7lrGNVjn0mc6tVLpjk6c5ZcJKdz6cONS81ObktjfbjQRywW+fPrnY9TpSLsxzuT59YOK/wBOPXvNtsRGHVjrL8+vm7ELvnduuJyzUnDncpz7dGb5beZvHoHXnuI5OTO7LjrAyeUYXv0crXvDiBO7HSaWiZec89ewevzyRrSo893JrPU8k83WJt9l9fk3LyFc5dLtucFnh/i9Vp9HD0rvxyK7i9k3M7zBx4T4PZ7H7fLbN82tIxq97YpUMXyrF917ZkAKxc2ia1VRMqaz7K33WcqQVlgNJ5Zy6cnLfrvp590UfGrP15dCcleOeT0z016R6OUhc+f89XXvxySNmvG/F67xrN2789pTcy59+TIDO/KvD6/SO3K0dJokit4sm8IqeN0zz9vRdJio652dOcvZiUbHSF47vbedaOnHs3zlKwTz7l23Rc8dq+nT05SWsS1nMvmfLpKWXPHavSTnXn1XPecS+b41ZdSyY60WS0deUinavAvnkdfDv6O1ydeNf1iZl583kSPsp/HrfOuJHeIipY483ikz1Khw7yu8Wfry5a7jkl54kFqnHtH3Nx78HW2uXGuKSxzpWcWnZ1e/R5+rRpzZ1D5XBuCjzLh29E9Xmld5VnNi17n0v3SRMeM+L1en+zyWHrjUR+bW+XT0HrnmTxDweu9+zy3DtzxI3NrXHrf+3PGvG/n+uX9HH0308NJyS1rnq8dGSea+bry9eXrfRynHFbubcuawbPl/O+8b1y1yxTZi4dJtXmzPDfF6vc/VxkNWPkoHLd/9PDoTcng/zvoei9uV574i8qDz1ePV5+mzrTyTw+3fz3637fPHY1RMW4ery9dnVZ574/ZW/J6vZ/d5SWiZzZvT55GzpSr8e3nfg9/pvfjP9JQ8yyejzzGsb7IfOvNPF7JcvnfFKzJ3vxsm8b15JaD5vRHculw68q3LN9uNx6Z2GuKTx6wHLrL1za5y/fjcNN0K2sct1bl15cay3znu/G52THPt28e/F05RSRCUDN7M6lKv3Tn1mKRy1iWuZpjpzHovfjOWKzSlQxqJzuamvPeer925XHphmFleTg497pz6+NYsp25ekejhsMErubDcu/ptvk/HVMxr2P3+KTsxqNyq/Hv6buVrM8F8Pt9h+h4bj15hpTzLzen1Ptz2XPiPi9Orc9l9vj2GFnm/m7+idZIXNRxfC/n+73z6fgndYCoc9zOlgXTc+EeT0Wbtz9T683HCVbUu0rKrHkvN730vYqTzJj0TQMLPDfL3sOOnrnq4NfMOW7r38/ZqYlT5dPHfl/S+h/qfPmVpvPfDvlau3JmlPEvl/Use+fsvs88fnVEzLt6fPkIpPn9Hm/z/AHe6e3x2HV80ytPo80hqBxS+UfP98zHsXfHn1z0dfPZumGKqhw7Ubyer0nrjPriPvKydMddZLxFC83o041K9OWknumLHvOSpKvz6Vjl026xa+mMEm9OmmckVDnuOy3azbM9MeXWvdOc9vNPzbe1bkVmqyDy875b6dLD15VHn19N6YmDGzQzSca8749bx1zz7xpx09N6c+isEipK2Q3PpP8u9b68bD0xb9Zzs0FP571HPw9FeZke3O39eU5Y7IPFgOXe5befcN07nv0P2eSx6k3ZhZ5r5+156FZ5R5O8Xnfqn0PBIrKXEDnUZy62rpILM8d+f7rB6/N6V6eHYd9xQue/RNWMWtc9eU+fp6J6eVw3nuOa5j9SbzrgWqYtLYvee1r3ntuaTcXOo1eYo/HdI8Xr9g9vnsG5nc0PC+duMTNabKB5fTWvH6/bfoeSSso3LVp9Pl3VHLqTzb53v1Y6e0+3y6pqpOd49HCPl4LMI86+f7njr6b7PLDpLdOM/vMQ1zJrim+P1xHL0ei+ryRlzcOvDp1YmXRYs6qfl9NY4d7b6fLLdMXPpjmWMswuXLS/L6qL5PTbvR5b735WbriJl4dZ3XOyWh+X1VDz97338959HHv0h15Ljv1ma49vNfH67f6fPZrUlf3jRLGcelV56pfDvbO/L0z08J4wqE1jiygOHeGma3y7y+p6l6/LNmuyBqMxqI5b6N86X5vV0V6v7fFJLqsgiD5dYvnbT1x5v4/ZoT1/6Hhkq03MIVrzd9q3HpnzPx+it46e0/U+bJGioaKb5PVbOuLnqeO+XtUOHf3D6vy5iuRYaaofk9HrHo5SLPj/l9FC8/f3n6nzpvU5YrudQXPfofRIs+Weft55x6e4+7yWGzhWnZvRvFtzruqlZvm3NfJ09H65jlo15dU1bN42WV3OvEvne2/dceverhwTXlXLVy9PCd1hpwL4V8n6dm3n3L3eWFzvyXz79H9/jlkLOSPGflfU3x7d7/LAx51x36f7/AA9xkaY8s+f9CueX0+x/R8EVN1TD1b2+PplaYVQPL6qJ4fd6X7PHX83HefT/AF+bauUYpUuPbzL5/vlN4fTjYvRx9D7ctgzCyv435r4PdDct9/fhfvV5rt1xtlVmuyLl8/8AH663x6ZdOXovo4XHrncvfy693Lvza567nVZVYoPOxGdzk16d6eEw1lGu502U7nvz7juOx062/U/X47TqZy6tZ1JS+XSAxvjzar5/T6j7vFeevPZNarnVc0bj1iMbtGs+NeD33P1+b1X2eTfLhZquaNw68mOnoPfh4l8/3R2Ont31fmStBpSicO3RN+obx5Nw35R4ff7X9b5Vt68840VQ/P2tWraLmvp87/L+ldPb4/YvZ5dkuCUfn0tWpOtaLnwbw+rm6Y929Xn75caqUklVgmklLjzyLNz6ep9csgdYhIteslmk8J8fqj/N6fpD6Pi7JYKykZX7vxDBKDw7eVfK+r7P9D5/ofbNRzahmei+rzsSRsvh3x/sSWuftv0vn1rHWv4ej+vy7ANaebeL3ef+H3ey/Q+fnvNe569B9Pl6qyrGq/z35J836Uz05W70+es8unovr80pqZwVyp5/5PXUOHS1duXXvnZuvOe2zCzWlf59PP8Ay9+O5lLLb2xaOmN47MTnsqPLdN47ysuGlyz0sE6V3pwoXDtjvG3fPiz09T3O6Vxp1NOs1TDznzd9m8TW5I6ej7zsy16mm5g5fMPP16Z05olOuLp15WcVmq5jzzXz9uDOuuagefS6+zy3PeJRddxqrz3z9thFY3X+HXp6Zvfs8to1OlNdlT5bicdJ3eaj5fTQfN2v/u8lz9PGwXCsj5fNvN39e65q+deV+L0wsewfR8cxczms42ed8t+pXUQtQ578t8naZ9PD1bvjviW1mpMzbUhEI1TOeoDfPg8vp9o9PPus23FEvO7VGrHr5/5+1S8ve3dJ6x6uUkz5NiejejhlZBZ268p+f7Yfzei/+zz3vvyp3OTfXlZu3PkiEl2XPkvyvq8vPd39nlsHXlDYej+vzbKiMbi9TOXyr5f0lnV29fl5Uvnp8s1uKWuTWGs8vPfnfg93Lz6GufoHs8l79HLcvBFfsk984fj2o3j9cB5+909nh9D9PGW0ylhSGuZneIXl0ovj9kfy6eje3w2/tnplVlYl5NYmdZhsXd5vXFeb0ed436B6vNfPRwkZrTFfWRzqX1ivSeW+X01/j6PQPX5PQu/Dua5VgkkZepnz3j08+8vr5ufX0D2+P0j1ebsiPWHllWYjGvPPP24efWB8/pvvu8Xp3t8W+WLmo/NkrPN/N3sfXnWPP3pXk9ly9nj9W9/h3zUNLomtWZSvP6L96eFF8noovk9Vr9fl9d+h4uiWBzvTJS/P3tfbnP2+feTt515fRbvZ5vZPb43NQed8slfzq+XUvc+Q+brTuerL6OftHo46ZYfO6zec41LLL3NCxaRm8HHr9Cerjz53ElB1xttspqdtzT+W/K/H6cePb6Q+l4+LPSjsR8ll7c53WcrK7z34v8r6XRL7P9PwZ15r5e119XmlOmJfWcUis68Y+R9bTjXr30/ncs1WOO7h7PPMb5yKKo/N8h+Z9KI4d/Rfd4YfOpnpym/TysOs9C4pxR5l4PbTfH7evfOw+nyWn08pvtymrNhiaEpXm9HnHz/oNm++3w9fbNn7cpWMjXZrSscuvmvzvo4s3z2+Hr7ZtWp1GCKzu5dqH4vbc/b4u/Ot+d5LruefeKYxQfL6Kr4/ffvV5vTPX5JNduds03PJvn5Z5+8Bx3WvH77R6fP6t7vDPbzuzXGjU4NTxnwetkP5/ThN+q/S+Zc+/DdnQabIyzxT5v0fUfX46N5fXUPL6rz7fF6r7vF0TWS6LiAjyj5/0Pavf4qhw7eU/N+hJ9+PuH1fmySZy89lL49K7y6+perzxnHr4P8AM+g+nP2f6PhtfXGyXTZ5t5u1r787pjppuPnHwevRrN99PL1Ttyzl12ebTN9blDFPPcXz3nrm5d/ob2ebtzrXZ45men9cbzGziTwP53u5OHf1/wB/k9J6Zhd48Y83X2P2eXcI1XPk3h91K8Psn+vP276nza/jXnnj9fsP0fn7wNVlb49fGvk/VM9PavrfIgMdIPl09a9/h2mRickvkXzfpU/xe2+e7wR1zPbx6d7fNnTRJqSnef0eS/K+r175Svfz230cPQvTwzsFxTVZHy+Z/P8AoV/nezrwv/o43XrnbSRWarNJT/N6Khy6a5PQPRwtPSb6Vkhx793Pro1lxo1nC5iJKFz1VefWzbXztxmbOjO8pdWpz3EDm+ccNxmenLz7Xn0ef0H08OvN3TWFnPrMPl5V5PTsK15vV17z7F9L5s/rO3OsbNFzFy+TeH23j1+ai+L2VTy+q++7xes+7xdGdM1azwyeReH23f1+btl8S+V9Naz7f9X5tl3jdLqrmZ8o8vpv3p89gm/GfB6qhx6znp4e6+/x9Mrl0az5dw6+nbTMtUTwL5/qmfTx9C7Y9E3jNdaecWejZ10mqzy3nutpx8evrffnb6R59vjMzU1qY2cB5B4/RXuPWWm/b/b5+3fPyjObGtr7c2YFX578d+d7+Lz+n1v6Pzu3tz0Zcmdeg+nz50k1J5z5fX5t836PdrHpP0fBE41ry9T9vk2GQl5Dybw++qeP1WTv5pnvx4M69V9nl7NMoVmuyHzrzHxeyC8/Wc7+fc16Z7fHL6ZylmCarK1y60rj0jsal+nGTz2ufp8srbmY1gmBROW4mMc6tGpw43aM2+Z9Ef14V+48s8/ftt2axYOuHrFhmp+azmsLnRrEIz4/4/Xpzvu3m59+Ej25yGNWJQ13OjUp3N5R4vb2zXHjfp/v8Uj259+U5YmdOpAY15P4/VjnWjn24Zr1f6Pzu7piYllqwueZnx/x+uyduVG8fs4ee+ZPX/p+Du1mYWQs03PnXn6z/XnHTVe8/ejeT0bOvH1n28JPUmrOvWYXKqy3mbj2vNvJ1rUzL9s+kdsd6zlzvufMrPT865ZYtql5zAJq57tjdz6pi4pe+OrOrhvMPNJfJPJ6IyYi/J7PSPb5bZ156+vGm8Ovq3p4iVzHSS3il8e3mPzPcTdk78fQvb46vy3d+3Ge641lZx0nenGoef0eV/M+jjNSHTnZvV5t9z6l7PJst5Mari2DpzgePbyb5n0OTn03ak36PL6r7fJNbzksVLCXNh3iJ59fLfn+3j59Vc+je75937TeZFcl4tYsGs8ebSfP6Kt5fTH8evovv+ffPRz7JQqhjvnPLpSAxug+H3ZeT1+6fQ8Pmsx5v4ffY+/L0X2+Owax1K1gzn57tdzx6zQed8x+f9GW6ZtHo8/oPq8/dZlmw6x+NWrWI+zznjugfP8Apdiyvbh6v9DxS+s5Sw8sfnVi3xq/Pfmfk9MH5fbus275+s/R+fa+3LZLDzXHnU/vl5F4/VLdcRvDtS/L6lc+ge7yel+vy7pqGzrkzerWPOPN2uHfEprHiXy/ochOejj7n7/H0TUPnfPJWsO3pMF9Fzr5v8Hp6O3Hs09h9PKcSDz01XNC1yuuO0wsrc+ZZzWJd2NzEvrnaUeWH1y50sLc1qddxQ+XTzfz9Y/h0ndX1D6Xg4cdKtytt6Z26ti3jJOdPD/n+2K8/dZ16n9Hw9e5QfL29Q9vl5Fs2+eZrufOvJ6/PPB7MZqb7c5Prw31dPX58rLDvLNaRON+SfN+hGceuEsz6fLf/V5+vpjf0xPWZRhWlKD4/XSPJ6+Hl2s/r+f6R7PNFLN9MS1OMbNaQmN0byeul+D32D1eL0b2eTj2n+nOUlEVJOQ2cO9A8Hv884d/TfoeH0H0efsNs1szptaLiI6cqNysD5vRSPD9K4+vy+j+zx2bpz2y7Jpy6bIjpz818vaO5dKd4PpTXXlcvX5fTPZ5Ok2ZrjTUP0x5T4vXy81b8f0JLfPPePXPpfPs3XjuzrKa1XMPvHjfzfoWHtxkjzfwe/LWbD6OPsf0fn9Eu3OtZB6x4j8z6Ppfu8Vw6Y818fqovk9WfTl6h7fPfvRw6M6UQNeR+Xt6X6eEvuZcOvz5873d/fz9Nvv/ALfL1yhUjyvlr1Tvi543hZ5RytD59N8Tk17t6ecFvFOkq2HsPSdBhc1mb8P+d7VGjj39s+v8ma6YrHPdJ8vo9q9vm3y43Omyqc+vjny/o443vr2v6vyqZy6wPn9Htv0vn74ZhZqs8r8HupHj9erG53vw6u3HDPT2n6Xz96YGw11x5eSfO+jXPL6ODHa7e/5mLXrvv8XaZWYmuzAheXTyf530at4/bbvpfItXo8/oHWdVrTG5xTVWpKjw7+WfM+pN+rwTe83Xvyse2VmKYWYp3cu1M83rmvR5ZjU3TWzOtk0k06zCMUjjuu8u0dz72Xvx9O9nk683bLnNC67nkuaBiVnz+iE83sjOfX1/6Xzrx34bJdkrjVZzaz5P5PRySwHm9cLw7ynfh7P9L5tj6c9s1nm4WaNZ8p8nqq/HrcPRw82+b9LPWZDry9x+n86V1NmazTZ5r5u9WzfT/V59eb4n8r6mNxLejl7x9Hw9cu3OlVM5ap1z6L0x2VSvL38t8npl/RwsfSey9+O2aIhLPK5PVtp7nvXqeZ4lQxvrWP56+hvRmO1mo651PM9duszCuW58O8fq43OI8vquvo5em+/xQON0rj19L6Ynt5LNdmlPIfJ6ql4/Tz8u9k78b99H51J8nqunblefRxyQMLnQeO/P+hTvF7Ned2z2eIWV6c/Wvd5NicS9SOzmPJPn/QpXi9cr389k9Pl1536r6/NI7zkJMa1pynmfh91P8/bu7eax9+HoHXM1pjZkJNdmFc0Ufh3qHDp3XNg1Lh35Tmrqucjv5dezHXl3zzmsprErLHZrFS56geXaPlwt9V9Pnl952Z1tlcuFkPrnX8arWbF8e8B5vT07z7D7/DP7zslzzQ0WcmseR+Xvk1Def0RnLq949X9/iu3bhszrJUc9x59w6+d8O187Yovi9vHm4XPpP0PH6R6PPvzrKXCyIZ8W8np9G9PGPzqr+T0Vbh33deFs7T1b2eSVXLNwryflbH1xjHHjrRfJ2i7iS6LJvPofWWZEUhirazb2rnjdJKRx6cO+fQtb4dPVu8uW+dL3zqWZ6q3J1rsr0151y3V+OuDl128+3o3v8OWpIdOcD5u/rPq4Mxsg5apy7eY+Lvo498ltPo4WP0+eo+fr7F7PJM7jRWaqp3Pt5t4PZC8OpFi78eGrR25er+vzbaSch02VXGoXl185+f7sUtXr8tb8/p9W+h825buaFYprqHlr2FR8nri8al/R5ezHbC49N9XCRpWYiOKSl43MaVDz9jF2tQuN+gevx3THWbz259YF4mfNcPPfJ67BqdfTHTvN97+d9OcRz63ZdkpGrWatefjPg92/PaY6cYPj29A9nlvfq81Zxq4L1S4mjWeK48i8vWA8n0JDWODGurpj1z6PhVzuxuw3KXRrFP53yjy+nPHXj4ejq3zwubT6uHq3s8ld5drhrGRo1nx3ydu7tz7ZvzX530MrzWsrU9g9vnlOmJPKS1OdPHeWrx0xA53XfL6Kp5+st6fNt1q09M+qdMR+d2C8/M9Z5NYsc3zc+ujrw8y8Psle3LIr3Ddu74l+mJPeIfXOy8+1usrs121WMvKvN1xl4PP3146+mfR8ElvNUw9Y7YlNSIlwWQufB/D64nj0ed451Yu/GxenzwXHftHt8vRZiU3PSx9OemPFfm/QjeXTGXnx0m/R5bV35eo+vz7KcVSJDeJNYHnvyP53v5s2S3mF49/SvpfJ9D7ToXIhIhdYs+plLSuHXz/yert6c4Ly+zt6+b0/3+G3auxeFKZLdOmN+dabKnz6V3j0gvL6q/w9HoPbz+w+nnv3zqTHnPHpRvD9C/erht6crb2427ryzXEiLIXn0vS81xQszyn5/wBCTupLeOLOvVPd4bJ15uVWVXO7RLvuYzXPyDx94fze/t1jjxvr6c/Xfo+KZ1zawk1rxqw65V2PGvH6pJYXzerfqK57umPbPo+DtNUtZ59bR05VfDyzz9fQ/Rms+brUPL6nrOW+cjrXvX0PBtWHzvbJX8oPeNuOtl7cPIfmfQjM2b9PnxavXbn6hqVQis2K6cN9vLz6THTlKTfjnj9El0xlqRHDpZOmbz6/NX+XXZ049Wdy+d8epdyFTxHzd8GIvzenHO7R34+g+3y1fGt3PV8789Dc/c67Kbz35F4u+OOizvCX1D3+Gr8+s3rn6b6uFNx0tXXn0zOFROdeK/N9/Nz3ic+Os96PLZ+3L1D18KtnUnvEsMwsi868j+d7onnuR1K9w9F8+j8j1T0Zjp0itc7TrO1UmJFy+X+L182NV/y+zv6+e6+3w3Trmr53du2OqGJMbOGKhy60bx+vR4fpeq/V+PEzNe49qV4/fZ/V57x6PPee/n6azlylya1pAdOdY46iOai+L6O2dJfpykenP1b2+KQsyayla6NYoEndl535e1d8f053rw5perpz9f8Af4pjWc4a66rtzVePSk+X0yu+UB5fZsV2LWfZPoeGx9OezOmvNc+fc+lD827R2zbOnPx75v0Aesaq9W9nC/d+G7Na0Zmhcddt16B34x+L478z6T3zmPRx3zXoHfj6HpEXFR1KVy11lp6SR1zk878R8fplemeZnk59JZPQ/d5Sao/LXPE90WnWbbz3o1PE+Oq1x66ee9fPomvafqfNh8dKHw3ce+PSdztTVZqs8T8XsgOOsc7xzrp1n1P6Hh8z8npsXfl6j6uHbIIqwqvc9+N/O92rGsV4uXaz+zxZNene7yWSzZCuUmFckvk3h9ta8/ZTcTx7XT6Xx7Z3zeus3xkirFMKxZovn7+f+P2Vzx++w+v59g9HmtfflcdupSzFMbEYVB5c/m9Uf5+0JZS+HpzX3D6fzJ3Wc5clzzrNQ0s0lzp/n7w3PtSvD9Gc68fR/d4vSfV5ck2TWc1koc+sVm8aB5vRQvnfVJZPpzkuvP2T6HgldYzjOUNVQ2s+EfL+lYe/mp3g+j0azu1l3Po3u8npHp8uyazmnGizyrzd6Xh6/wCzh5h8/wBsBw756xs3ja39CfT+Z2tb86ZSt8vJfJ6Ln35XLead5+3mng92/rx6+uJCz030cr5UJrnB2edctOz0TpMtY7M68O8Pt7enLQmvl2kF9Q+j4M82r51QvL39M9XGZ3m48+mNnknLXnvn77M3Rz7asavXs8tq9fl8483aZnT1D1eadl12a7IHOvDvB7NPPazrmzuw9uMt6vNUPF7vevp/Mmt4diMbMKqfHt5D8726c6j+Hp7OvK4+3w83H0e2+/w7tRpjZimNmhfKvF66D4Pdyc+1r+j8rv6cfQu2Lbqqx0rMU1pjUHjXjvzPq87Hb2881czPXleOuZm0sxrBCsU7eXbzHwe6tdOdz7cbt24dNuc1lLnK2sojXPzvKI4d4udObG4Tl09i+j8+7deTXOXOacuNiuai50Th6OLj6Kv5vTzRZ/R5/Z/oeKRudkuUrMDlufDvF6mnHy7wfDvt1np3iy+nh7L7fFul2TWUuJEs+BeL1+l+vzx2L5p836W7eN2+e7eb92x6l6vLvzrZLxWeOcro1LV1z0s0jw+yq8esl34bLqwdefqPTFnzur9eFQzYK472+hLHrMvnp4X5uk50kcyufTi5dPWPo+LizrizuGZ7sdJzryuWdSDVNk8f8vd6xwcO2rO3np7B9T5sfy7Ujjq+enjf7OytdmrWfJ/L6Kbw66eeuPHbTjfpv0Pn1/G3nXtvu8e2xisxMKoXDr5N873aMdd+udq9Xm7OnPZnfr/p47LHYrMEwNVebeX0+beD29vTlK9/P1b53LpzvfSuxhZimNarnSUHzeig+X079c5zeOqrV15XDo21ijsRI8+/mPl9N19HlltZBrlKTUYhUO50bh1eO3EsVy69PTn697fJJ3G2a3SuaxNVlYZ5WKbx78vLvDcO2ux9OftPt8kzvOebsgXFNOs+T8dxudHHtXeHpVmlnt649i9vksu+eyaylF0M+HeXro3n0rvjy75/thOXU1nq7cdPPt7P7/Jdt8uvHQjz7fKgct2vrjZNcdx578/38tzN9ufLnc50xe+uL/nVF6cOBayzMNS2pBTMhz7+d8OkvuR+uezn0hOW/R/b5ebO7LvMBrljx9Mn05Tllsz08ixarx3HxqzebHTTy63D1eezd+dYwsVsv25WuJeuFKVnp5J4vQZunOs5eiz0T2+Sm41ctPSfRwyoMbFVZ56oPn71Hy9tq6pbJ6PPnp2b5+vd8bbGJMaxISWnculF8fp5cWa9HCW68u5dWOtp9HkuOtJMaDXWuShcukfm1zl0lt52ZvfrKnWPvL1P0cpJru5dqFi3Hpz6hq5py1e8/I+HTTx9Nm68dzUJjcdz6ekezySPfz9Od2CzPOtkrt5rjy3PPzH5v1/Rvb4Y7n1huPV2S3Xn637PLVMavW8bZSMa0azSXPy7w+5cfR0JspazhrHrfs8ysnbmQVy67PNsTzzz9pjpmu+H6HTvlhc4659vbHRz7+1e3yasbs1lOuY3WaHztx0h8684+b9Hd04dHXjYu/OG5dZzcsvblG41Z+vNFUYmW++yp8t8nLpB51LdMcWsbeXav8quPq9O+n8zsm8OnKK49bN0zp1iE5dJntypfl9VY5XqsjuXXXjazu8+zySm5AYvofo5LWbxm+e516DvPi3m703j01c95TSl0Z1Kd+G3pj1T0cLf1w7GREscWPU8c8XrqPm7Yy4yy/blE8PT6L9L5PqHRsrJGcZTJq77xCY1474PZGc9yXblYvR5qz4/bjZ6Z7/n3jV3UjWlBxu5deXdNVXnvzDy+iT6c+6ys+X1ac9JL1eH0TvxuWO2y3znN9N03S6E87mPNvP2jPN7bz34Z6lf5de/ePVfb45rULKhlY87llSctz5fnHmPzvq331cIfluM57Enu/P2P2eTts4rKty63rWMTTrNYvLx75/0I/z+vu1h2OzHWfQPVw9P7+bVZRuXW97zmkXqeHeXpvmoDye3r1nKzG56O3Lg59PZPZ5rvrPlaXvO4zpirYnFZ1Y69Vz5t4fY9c5XvykumOXG7L0zP9ecTEfy62Lrzrd5TM6wXPpPdeMBx3G53L7xB3Mjnde5WN5dvYPoeSu8O8t15REtlqv5bt4ldTk5dfPOG5PpmI5Xl57WOk11xd++KdnNx3qW6c4bnrh7cPVMdeavnvx+nPLDOsc3XNcWNz3fhnqe1+zzyOs6SoZ1dt5E568Y8Xqr/n665cSX64rXm9fq31fi+la3upHnedXbry6pSIyzx/w+2vefr27xO+jhUPF75Dr5/QPZ4vQ+jqqi51K9eU/LslRx2eXeb0V/l0l+nOv+T2QnLpePd86057en9+dZ6cq/y7W5jzTOYHl0pXh+n6T6vPv3zjefSzejh6J6fN0SgzVqUnFvc3oZ8sxnzzw/QtPbHeRWNYkz25es+vzdMZNa6gpnkx0s++cFrj4l4PbBeP6Vi7+doWY2T3fj7T6vK1Zyp53z6+kdOXmPK0Ph3786huHq2ayXJrHX154Y6/RXu8WmWi7xW+PW6dOdH53Yt6658+8neoeb0vWZLtz26zsmpjcu/p8mqarvPW45evLdy69OpL7xUOHaucushvPJcbsdY3F4OPT1v6Ph77ahx659eMxNwyWXpgudXHv5v5+2u4Wd8XLamsY9l+j4aRw9DuLh250/K09edlm7ly7+V5eX8d5c94mObrl5c7snq8s7p6v6/N5bz36j0x1riirhjxbxeqL5bwlxO/Suce3rv1Pjei3tRJbP25SudZRjWCc9eU+T0VLz9urWZrrxo3z/AKlm9fgtHo8850ytW4bzvjJcjFFZUueqBw7dms0b5/0995X7ry9q9OIjrw87zmF5dOXHSmeT29l1YO3Hizr072eO69uO6VrlGKhH750HEi+PSpeb1RHD2Wbtw5M6xssHfl696/J2mUuSqI/WfI8SzWUfjaR837Vn7cNly7FZu6Y9x9nk7tYzmtmdQOs+f3Mbx6Vrjuf6Zrfj9u/WckWp0dOcRz6esevzekbzW7mGqNSkefoaxbt7tnXj5F8/2cWdZ752D0coTl0tHbnO12deWc3hm0Llvf24Lj3vXfllZVeOojO5DeIHMmbqNxqF49PRfVwsHSV3j1rWuXLx7Xv08um5LMlpnDrVePSd6Yh+OtWd686tvo43rvjyXy9ujWbn6eMjZss9F5d8Ln518vo54xzSXXLplwmpr0+Rzdh9njvN1aJpIqxSJl8R8Pr4ee8ZWR3Lvt6cb/8AQ+bs3fU9ztzoTXZjWKa08x8vp888nqysM7iuPou3u+ZNdedo7crZq71YkEa41GR5Z5vRWfN6K35PdbbPoP6nyvNHKN59dWdV7l2qPk99v9HnsHfh6v7PFIWZKzZNbJVLquazcUDhuN59aH4fpSO8zu+RZY/Ry9Z9fk6DKVrlLrSr3NPuIPhaP4Pq6OXaw9uG3USLefYvb47Xvm12S6YqOkTJ5F8/2z3q8kf5PZHcu+7WHYazt6c+Xn2+mfpfPkM2j7wprhPL/H3fTj6D35yK+MfL+oWPWNvTlzY6dm5bevO6+zx7s6051QePSIvOZtvHbn0alL8vpo/m9GWueXTlnjtq571Y36D7fHaPTwrHLdVmMuHquvq88tvOy512eb+D3Vzh3k+3Hm49dcqlF9a+l8yhcekT5/V6B7fJIax2azPtXDn1pEvhXk9G/Nxl051x46cnPtcff8uG597d34XT0+e02y0Y2YmNQGb4f4PXpzrXnUTw9O3ebr9P48rrNy10t5sTGzCzExrBmicPR5h4vVE8e/Hz7XX6XyO2WV1LB25Xa3oosSKnKjRrNA49fHfmfVmuXb0f6Hy4tCbr+WrPWp+b0+j+7w+uevydZkuUuS7c6ZilIYpXDrozuLm6j5PZtSR6c7b6OPsfr8nSZrlK45Fp1zB5sc5xXL0VXx+yN59Zbrx69TO5v3q8/qffztc83KWnakBLSfL3qXLpbOvGk+H6Xf149u+WzeOzry4+fa+d+Xr/AG5RSU44s65U868vfv3j0j2earebvUvL6tmuff25SnTEJz3dPRym7OC4WegsJx6cvfzymOnRvmazwcekdnfZvMQzYLrhyrvDpY+mLF6MSM3QuVyzqzdufJcZ3OWpv59Khy2132QvHWjO+Pl2u3p49elG469F746unPjuM9Ztmd3Ka8G8/aFTRz1rzrjx04eXolO/l9D93g848P0fQ/b5O/eL0ky1jZjZrsqeb474vTyY1F8PXu1yuvt8XAxauuZu7slk5YVimNYJhZT+e/FPm/R0Y1Oeny9/bjI5sjUn053nclLoRWYDMLNaRM1B+T2cvPXHvFezrgx01r6V6/Jd+vHc0Qxy5KRDpTs5r3LrvbiM75ufSMzrkkvHp4evenz9BlLlLF1WTnXoiBcorn24+XWucO/JHdvEjrMx35+0+jz5mzNiVrUcK5nknl3N9eWrj6a/x74syHXl09OXb0zAeb1/R30PFySVc2ze9YjCmOdkurl25eQfP9sdjW3eJPty6dTjix9M2TedlnRnamqrhj34S+OsnrOrWarw6QXPp06zGXEpnrpiA5bmt59Q9nn246U9njxbTtnqK412cvPdJ8/eIzrvsjOW+fG+fn1k+mPW/oeCm898vLrfPTxVxlTublnal+cvH6s45cb5MdMJd2udp9HCQ7+eH4en0f1cObWOlL210mFzhXn3Hp414PZrz02XO7UmvRw7N8LX15TrrpssWszkuuxGNmmyt41454fZH8+m3fOf7cpneN+ddes2jrztrTpIlyEiWQ5dvPeHapJDY32anrXr8krZkYhDXFRIFKLznHy77WoqajOXUzpWWLvw9h9Xl2rsla88VmuaMlhXKC59Yrl2huHdRprZvHZvHuXr809ckvFFO1d0qjzfjrl3zmc6p/j92Bpud3Tn17xpx0s/XHuvo40rfN52S6loXC7O/GyLJa5+J/M+plc7dZk+uC5bUpuXHt5+zU6s6wap3O9XfhNY6dWsxckBy6QWOnVqcNx3Z6EsHhtPSfX55uapebx3Fvaz1FrEdHRLVePap8tT3TMXz3Hc9acdNh6R7fHzWwuV1uu7pgZLOvUuPPr4Zw7V/M1ZvHje4zMmbr6vPxazKblibVzI2XDOsbMa508P8/Ws+fttMJdlzYu/LPXOx9ec+61tj0W6kRGNmuzEi08h8voh+PTK5m+uJ3pjVz6dNTnXjMtwdx6A3kJNk128+vg3k9Veubv6fPN753jeRcZGuUutPJ3KC83ukd8d2N624XHSI5dHLnqeiezyd28X7WMjOXnKwmpaVedM8H0LX6fNy4617z93LlZjZlvn6d7PLLTV6ucIp2nOa5YLDz7m5OHq7zTKWa9Z3dOUl0xVfH7PSfb5Oiyx9uezO1Lok8155sHSV7nuC8fu6d8st8+zrib3mExZ3pO+zGXTm3brnCWnTPb25zeN6krGNVTzem0ejz9OpBOcnnrsWCzmN56751tvXBrHJ05z2OnVvOGs0nhuVuubOoSZ3aiiC5Ux0zl5sdZvty6+3GTzu49catZLC5q3Lcr25+a+D3dW+PLz6bDKXXHRvG7Pbl1y9O9vl7W8bmxLYM3XZR8dLdvHjHm7VzlpS6o2alh78dusQPj+j39/JcPZ477nrKNa0ViSgc+tz68qXw7eZ+frpiV64tHbjr5ddc1T/N6unrw9B9nk9GnTszpWdeOvh/l9V+9fhsXTFLSyZ3I2Eua8bPljl594fe+fe/eny891F89xvPo5crPUPb5bv05VizoxuyWYRVdTTLB64eV+D39mets9PngOHXVneVjQ3m7+nh6vvFIifl02QdLN0nnHLUTy3o4enu6c87C5Ws9Xbly8+m5r1D2eSnc9WJqU1Nc1E5zVLy5+XoM6huHfdvmb5yvXMtrNT56uPXHUTXXFT56s81321Bz6emZ/O6pz1Z+3HzfzeiX3ndcxVxJTruiJkhuWpTSY271x78NnDtL9cROZGS2rrip8O/CzA89TXTEHy1q59CaxzeTn6bj7vn6y+bbN4RGpXM5uXZX/ADd6Bw67pdeWSqMJe7piN4+q0+z519742Wu5t8sTFcX0yb4zwbzdYjGteWmXPUtfo88Ly66OPp3ejx+h+vzXWblJrGyCljNZuU04puN+Q+X0R+L39MWr0effnURx71jh6JT0eO8ejj6JbMTp146cNxr3zKLPPM30I2TUaz5czUPP1rni+n6f6/H09MRfLrGY6EuVz6Z7PLdN82vPrPkvLfq2pDVzEVeXm/n6VrxfT9M9/hg+HXlxvZY6dzK9se3duPRL5504Unh3v3SBhLXMyoYQ3k98jvkkysx1l7x19MVny+r1n2+WS68+eKn5+1+7YUtCxnZ057eXeG5bjOXU1nLpiW6c+rUrvPdu646FsnbjxXNY83ovPSU5z6Nzt59OQmuvLzDx+rs3NlzyXHVNdk3wRFc7vl9J9nlrfn9Mn6vLx8e9l6c6Py1ce/LdVc8/ph4rfNN7RvO82NmdYGEtm78NW5PtWvty1WUHjbh6eMjNa7PLPn+/Vcauewa4mCSe81jzev1n63xLG7PU23PnXDVl9HL07j6O+ahrPCPL3jca1xql3aza/TwqPl9Udy7Xn3/LuffncZvrs8lxr1rrnu59CMNZgJfHPN3guPTs6ZsHbj22U/xe2E59PRPd8+X2uu8W7l33rw9OWi56m6fvjXOPa275+d4RWNUTw/RuHTNt9XlguPfg56xXZp6b6vLc+nPOVJUdSpyw3LfovXnxs0bnPPPn/Uunp4ZHDz3sHZlZv6Z9q78bBFa6c6ZrMPi48+1x3nTnXmnORPDt0TasYrDWd/TnzY2l9d9fmLNMtfjXz3aumfMsc+nPa69efl/h9jUuejpiT6Z13MbjVi6O+yy9/NpWE56y59eXrw32w/DrevRy1M+ZeP2d2ps1Oe88munO9ERGLz5vrHt8lf499fTlnL2xH6ln6YyODn1qPLrA85Jdca8dI/ncM6U1rjNq8e3xRudXjaEkjdc7XudFZEXz35R4/XI6zz4uUuKYzW3U5OXff283rHv8Ei607lri6cbLqys1f+fXcVo8N83bhxpGrN7OmJzty88+b9Wd9PhuHq8lq78qzz6buvL0N0tHPowjVrMdrPkvDrUPP26NYn+uc7PNfmfWsfp8N378u7cnc69QnXl3zjd8YrWabrMDyb875MbqfHtXvN7vWvofPhOHfjxpmWnqPq8tz6c85XLWLmBOOqTy1O6xkxSvL64Xze24+ryx/PeQU7Nup6j6OHotnDc+f9OeE1xM0jj0uerDZkBhX/H9CV68skdK5z3jp3is+b0+nezz2ftwylxmoy5o3Hc7rNavOwY9Elcee+T15oaz1dcd+88EbyY2sGuch15ZrpPP/N2ku/CP59J+y3dc8UnmXk9UhubLOW5zs7c70kNhyY16d6vPunSgcdzXo80T5+939PHtrKzKKRw9MdMx0k1rUTz1z4YS65cJq5+nzRU1O21rMvHp5SFm4zsLnzzxeyGZeOmMIxlxNi17y+2/fT+Jce+POfN6bp6eMjL1EoXzl316zT08R83fnxojEk+meDl2r3m9Nz9/zJ/ry2deUvq9jVnls2OiEYazy3PmPPXn3l9G25nuuan5/TB+f03v2fPtO1g59fVdXm3ir9ONeuYVy4uXbVNwnPVD8nvsXTEvvGnOkm7U9Q9fkue8ZzWUtcuYgxl4aidcuXEg+Pah+H6U51xIa5sdZVnrNv7cvZd41WUHpx5ppzXLEFrnQPD7J/0eas+L6ElXRrOVjZN56umIvlvim/bfZ5C5zmsV5qrDn534vVPejz+i9ZUvN2rfHu9Zy3iS68+3ear5+0/159ult6c+jeNkqlqWFc571Z3e+/Gf6Z4pPNvL6u7ed+s8knHEpdYRG5vJz1f/AE8Otavy68PThz8PTdPT5unU1my54uXeNko/DraeuOTOuTGsJdUYZ10VavV5YLl121du/HdZhZjYWKPJPnfSsPbz8udY5qMDGITze7p6+f0T6Hy4+dbFq9g7lXEzNzk1LLS5PIfP3wzcJEvXqU/wfTlvR4rf6vHKbS/bjIN5k5FmztmS4Wc+sUTN8r8fqyNOelV8ntsvr8Nz7cLNjr7VO8brnVevKNc4XGjG+aagOXSmeb2ynXluZ0zWq24ejz+2eny5S5zWmSp083KXns4t8a9y61/l1qfk9zsxmiwBQ+i/pfOt0kH05VTUzmjNwmoS8vMPnfSvHt+bQPn/AF3NJRBFaJIdeHNz7+9/U+VzyZTWNnOsIz5t4fZfPd4dTNV+f9WH5dmhIbqrr3503nZ6N6/HPejz65eXNpPO80nHz9Ge+Np9HCwTfn3j9u/XPLXPlTXUjOjzrGFlO+nz1TG5azm6cYrxe7q78ereJ/eN9dOOkHJW+PSc685DPTnTKa1px5tW83t9E+j8uqctnH1T3p8sbZ03Mhc9eplVb8Xvw1xlKWbnLhcReNVTy/S3b5XX6Hye671zpyM6LnVcazv6Y9Wx3nD5+8vq4ed2amVzy89w3D2S/p8E924S+td2ub6Ywzrdq91z2XN359hcbObXPxvj3gPP0hOHq047SHp8V568LPnt/8QAMhAAAQUAAgIBBAAFAwQDAQAAAwABAgQFERITFAYQFSEiICMkMTMyQHAWMDQ1JUFQYP/aAAgBAQABBQIhZ+TzEXmIvMReci85F5yLzkXnIvOReci9gi9gi9gi85F5yL2CJzkXsEXsEXnIvYIvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZMvZKvZKvZKvZMvZKvZMvaMvaMvZMvZKvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvaMvZMvZMvZMvZMvZMvZKvZMvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvZKvYKvZKvZKvYKvYKvYKvYKvYKvYKvYKvYKvYKvYIvYKvYIvORewReci85F5yLzkXnIvOReYi800X/J/xAX/J/wAQF/yf8QF/y/8AEBf8v/EBf8v/ABAX/J/32ZP/AG/4PL/k/wC+yf8At/weX/J/32T/APCBf8n/AH2T/wDCBf8AJ/3uEyf/AIQL/k/7rfV/+ECf5P8AYS/4QJ/k/wC+yl/wgX/J/wB9nTp/+Dyf5P8AvcKLLhTb/g8v+T/vN9Z/8Hl/yf7BlL/g8n+T/YN/wgT/ACf7GTf8Hk/yf99vo7J/+Dif5P8AYcr/AOn/AODif5P9iyl/wcT/ACf7HlOn/wCDSf5P9m7f8Gk/yf7Fvo64T/8ABZP8n+yb6v8A3/4KJ/k/2Ufq/wDf/gon+T/ZN/B1T/8ABJP9f+yb+GUf/wBJyRZezBe43Mrku0jk5nJ1Is4J7JIs1t+I3IuzWRumJF//AOMn/r/2vP1k3/5bkjFPaGy95nUr0k9ifHaU357PKXRo/q0H5XPJSP8AiX5aEuYxfrJ/1d/ymdpJiPBewSKjckmvflrY0x4Ouef/AOFn/r/2zJlL/wDFkaEU94TJ77J783UrU085TXLMuF2eS/EEzO6lJ5P+IRh+XI/0h+ZF/wBCb9STbs0Z9o/43k3KaXK/MF+Jrsvyy5aT89UxpprhIprsl78OWtidRnGX/wC/P/X/ALZvo6duP99I0IKV8MVLRZPoEdPZK6eTzXVmTOn4Zcu6/EF+ZLs0F15Tz/MY8KUnk7R6tz5Zof7yd+GD/jO/8pv7G/X6P/Ln/dRl43lHsoz4d4/lp8v1eK5aS/aK5aa/Zk3Drl2X4df2TEdNaNFRvzTX2TXhKJxyXPP/AOxP/X/tm+jqX5/2/KkccFLRBFPpMpXyupWjST9pJukV+XXMV+XX6xX7Ov1guZSX6jXZ5pmjBd3IoxaC8nd4s0GkTtKLNBizdQj0iefEYs0Ynl1FFusS/kQn5GRu8AT7DmzTiInLTZpsMvEpM02YnjeTNNvI4k/WbdpDXMStzKC7QKv2iu8Zr8snnF1+WTzZMnkv1kvzFQtTZNeNFR1VHSE6jbDJNJn/AP0p/wCv/bN9OFJv9lOwOClp12UtNPfPJTsndftJeJk3Vfs6fqy5k6eLJnXj5XaMVxKS/Ua5lJNBorydkw2UytFNDsndot+x0zcMSbylCDDiUjCgGHH0g/lOrH5dT/013/kIb9Dqx/Llzyij8jBL3UotNu7gfldXGoFYjSH+WL1UotJdpwTPArdZRXkZeNd3iuITX7Mu0XXDsnkm4dcuuYrhfhlAs2TW7EVHVmybTgo6AJKJoT//ADJ/6/8AbsyZkT/uTsiGpateKfXZPpHkpW7Dp+xEwWZfoy7O6dl2iy/Z0/SK7u668rtGK4lJdIxXk5XTsnlEbczmowaKkVmfxvNfiLeRyKEGgiEYbNByOiFd5DGwo88IT+zNWS+IQYeIaf8Aa2nVR/6dWf5ZE/5YL+KaMN3cJmNB+JM8nqppM7TG0ngbh3/ZukhqBWmpDaS7TGmeJG6PFeXhdYyX7xXki68a7Siv0muHZd0zRkv2Zdorhfsv1XV08WUZcJj2IptA8VDXZR0guo3AzTSZ/wD8Wf8Ar/27fSbcp24/hkccFPTrxUtdlLTsSU7diadiEXrxTdYrmTrhdor9nTxZdmX7OnaMV5OV1k6/WC7ykvHynlEbd5TXjUiNBczmojaKmVoLiZFGLQaZWgvG8/oQ3DjF1dEM8piGwo8osnslb8Mmfz2/pWfsX6UX/kKxDyhrF8wFbG8oiKxRo0ZBnArEj/dO0qrxm04zi049p1lEjTYkGIu5AqMu7SF2XkmJNJps415ZQTPEjePheV4r9St0dl5Hiv0Iusory8L9JriTLumaElxJl2TNF1xJk7pmi68S6cKJCRdr1qCjqkZNrjUdKvNRNCf+/n/r/wBsyZdlOwKCNr1oqW1BS2CuvcuETxlJdBRTOuHdP0Zdl+XT9GXdfs6fpFeXlftJdYxXmZftJNGEU5mTRnJRhGKkaMV+81EcYqZYwXMyKI4wUyRg3aZVCEYJ5NFu8jqA4jZSLI0hiiJkUzykEUQxVo/RAEwBqybwBrD8IeVKXWND8VfpSf8AT6VX8Z/o39La+k/6KbPyynCYJDKxYKYZjcNhi/SQHZ4WfypA/PmmNM/ZnDy/co1AjEUhM6/mwUTNJ3E0l1JFeVmTjjNdZxXldlxAi6SZd5MuYEXR2XM2Tyg66L92TyZNGLriTLtwpMMi9ZmUWKNRu2IKOoZk2wyjrV5KNwM0zs/+4n/r/wBnOwOCnq1oKW3Dl9axJPctzUu00wWXjXEIryL9nXVl5IsuZuuq7wgvJJ1w7r9YLzO64nJNCMU52ZdiSXjZSJGC7TmvFyvxFvPyukpqMWgpmiNckIoQjBPLheeRVATRflFsNB2E83U5tCP721FmiyOeTzAFgQRjMAdSEn+sv6m79NCfWrCPWP0p/iS4VhvFa+loHnFVN5hqUezD5pE+hQzhIJomijV2KoHkN1MbTboWuhGiZuFKv1drDwTPypiaa/mDUCwIpDaa8UoLzdU3Em8DLkkFEsZJxRkuk4ry8L9SN4uF2JFMWLrxRXEmXkdl+hF0dl2my8kV0iv2ZeR2XI5Lqn5TxGmgyiQ8FHQsxTa8mUNgLqOjXkomhP8A2U/9f/c5U7AxqevVgn2oOn0rE1I9qSeE5r14Mv0iuXXEnXEWXkZczddOU84DXld1+XXWDLzRXabrryu0Brzcr9pJoxipHjFeScl05XMYt52ddJzUBwgpEjFvM814uV+GU7EBrkhVCEBrspWW5YPd+WUpxg3lnYQhQCyMeIWiJzv+FyrFh3kAEa8Vyo/15/pZPGuGkJxB+lx+5+VyuVUf+p+l4flrVjMcH0s/0lj6FHE0K5XET6Hrv2r2mN9JRabcEqIRoGii14kfzzrqMmkz8OnB0TWerqYozXBBqFmMn/upV4rsQagaM1KLSXjeK8s4KJYkTiZ1xOK8zsmkxG8a/mxXscL9SLxuy5JFeZl0Z11ky7EZeWLrxribLvNl3hJ+i/mMvJJl5IyTjjJSrNy3mGo3rcVDWsxUduKhrVpqFkU1z/25/wCv+LnhTtCGp7FWKluRUtazNTt3pu7TIo1YqAXXjZk048O8nXWTrrGK8rLmbrpJ1+ILycr+Y68XK/UbeXlcEkvGnJ0XllJdCSTD6qRei8pJLxTkox6KRuiZykTV03LKZei5MRRBw/5UzMNcGKhiYa/KLYYb+MxlGHRvyjWfG8a8yv8AlflHsvCQa7xf8r8qzYm0q9f14flflWySMQcGFD6WP6m4ufp/r1PqB+ND6OqD+Iv0KOJh0yPB+fpZDGxCraeT8s65ZWK7FVe33lyy/CLX/YNtpS/C/Cev4nHbjKX4Uoxk3hcKjbhzyynCBIsKQk1uLPyzogxlXSY17UYppRdpDHN+soL2YxTShJpCHJdZRXnaKjOE2cI1xOK8/VRKMi8UFxJl5eE0xkXigusmXfhdxzXjiuJMu7svIOS8cV1dl2dl3g66RddHXThPAbqLOyazbgoatyKbddlDcA6hpViKJIz/AIZ/63dmU7YRom1VgpfIIupa1qalYtkTilNPWCzt0X5ddF1HFeWC7O6Zl1hFeaDKU3ddeV44MnJCK7u668poQZOWEV5HkujyTDHFSJCK83ZdXkmHBk8oxXnZ11lJRHCKd4svMzrwymoBHBfqpGGy6SIoBGNcRRDCGuJmQxDEv1RCDFHtOwhhGFfhSnGLeaVpBAMDfqv1RLDmmAA68eWXLK1b6vWBGvHll2ZXLTVhUq/gH+F+EQkRwzYcj/C6xX4VL97H1h+NX62v6fQ+ugOUUIjGh9LdZzNUs+eP0s12sRBak0+foYETxYxKijLs3Log2LH+fWQjseP5Uod28RAodtpP+VJuy9eQ17MhqMuzccp6vC7lghl7t+U9blfzxprDc/lSC0l1NBew8VGfdpCaa8RIruSKYrSUh914JMuSxXmXHdvCuCxXlkyacZrwsuhGXYjLysvHF145Mv5rLyLiE14V1Iy5kv1devCS9JmeLWBqNy7BNsHgvvLq5btTtOCRE1MaYI2XYcF3X7Oui/lwXmiu83XDuuIxTniy8knX7uurLyxgnNyuSOujLlop7EV3JJdOU3EVI0YLzSkuJyUYtFPPhPa5XJppoMy7Op2GgmkYiYCb8J58L2XkvHOai3Ruzotphr+edDEwly6lPqz2iGQ6/V+XXLo1rxJq5Dv+V+VKfSPkLoIY/DDmS5dWrchvVrOBv2X7qc3hGrGdw37L9l+y0ZSPNuYt+y/ZEm8IZLS9L9l+y/ZTd46/7L9l+y0QSsVKZ5Wa37L9k/ZCeVG5zJfsv2VoBO1Wz7QuHX5R67WIQMStP8riSdn4esWsgWGsN+y4dFqtOXnJXUf2bxolaJY+uauh2oklw7rqvUZn8pQoRYmbhErxIvGUaawzPxynG0m9XouSQUZwI/VSrQk/jJBebooyjNnHGS9fhfzYprEF+HTgg68coru8VEg5JxwkvCzL94rysyaQ5rwjXj4XLsvMNdREXiguHZd+F5QuvGJ10Zf2XkgyaYpLxjVov9T3m6/mOujLs0F512K66SdNDqnN1Xlm6/muvGuereddyyXSbqEOqkTq3nd1/OkvEvyykdoLykkvGSSjDou0lKyuTzXgX5ZPLq3mlNeAs1ALDX5UysJeUpE1Z3X5X7IlhhrqcyGBhL8r8qVt5SapIj8Ovypz6N5jWkGt4G/ZfsrFlq0I1y3H4dflflWrUoSq0/Xbh1w6/KL20bDR4bh1w6m/SOZCRn4dcOuHWxNx0AC8YeHXDrh1abjV4XVdV1Wb/KL1XV11WhT9kFI/tA4XVdVZE9QopRLDquqIGJYNOefPjlcLhHpsVx2XHPqui6s6eo4nFaaUuFwi14Gj4i10KwMr9WXVkSmKb/zgIRhGXDJ4RknqtFeWYkIojNxFTCMi9d4Ly9FCQiN1ip1gzXjmNexGKhIRGeI3b1hL94L2oRUCCmpQHJeCDLmUV7A2TSHJSGKS8bMu0or2RsmIOacYnXXheSUU1ka7jm3jGuHZeSTL2RrsMi6DVsnWz5nX86S8UnTQ6py9V5punczrxum5inN1XlI64K68Sblk5+q8xJLgkkw2ZP2ZTP1XlNJeIklGHRcyU7HRdzzXrykujs37MpWOrs1gijVZlxJfsp2Wg/8AUGQ67DX7L9kSz436WDIYWEuJL8o1thy9c1lQH448SX5R7fieNQhX6uuJL8qzbccgU3afDrh1w6t2ZQerT9durrh1w6vnmyrVGqh6uurrq61HcrwF0j1XVdVox8lnquq6rqrzcaPVdF0XVWW9bU6rquqeKsQ+33uF1XVl0aTPH7WVuHXRl0Tgi8XjLMeHWcei6siV4FjwSghTGaHVl44ooBlj0LUQCisR6sujItYZm8ZayCYJ10iurItURl4ygQrAiP1iurIlQRF4yiUbQueIrhlOsKa8ZRr2oRTdZL8KdcU36EGvaaCgQZG/VSrimvHOC9h4IZxEX4ThE66SivNKKjYFJcxThE66PFeWUU1ofPaDqQxuuvC8k4r2oJiQkngJ10irLcWXJ1Xnd1yV143dNHqnn1XnXJpLxSdNHquXZPYXY0l4pOow6LmSc/VNI0lIM5qI/Gv2UzMNeYs14CzUB+NfspT6t5SEXqkmoC8TfsneTKVp3fwmKhh8Tfsv2RLXjl47B0MLBb9l+yPZau3Fq2g1mBHiS/ZEn44+WxcQKrV48SXEl+yJaLYnWp+tHiS4kv2Vu3IcqlP1m4dcOuHVyy1QNCoSK4dcOurqXLNnRe0fq66uurrq6ZnNt9XXR10ddHWpHra6roui6rXruWjVI1iv1XRdFaqRtAziSePDMui6KYYkiGT55uvK6LovGpgnnSFKBx+NeNOJnRaDjlXPA79GXjZdEfPgZ4n9d2HF28UV4Yo2eEyeJ6qAUVlujLoyJVEZvVIBQsC7dIrpFTDCcfT6LyOJDcRW8cU44unoD54MJQOGT9Ipxsp0xTfwlGvYaCg4iN44qdUZF6zwXcg1CwGT8MpChNvWZlwWC9iMVGUJrqzr1hrxzivJKKicbr8J643XheK6kVpubTdIruye1Bn883XE5JoQZdlIzQXtcrsWS6RTTZl5VK7CL+Ys105UHjBMVEsRgvcea4LNQhEa7ryKVtueDkUK8YLsuzqZ2G3tkKvXlNM/Vuzru6LfaMulg6HBgx7Ouzoh/FH2bFtAqsF+0l2ku0kfQ6ThUmSXLrtJdpIhvHB5G0kIfhhzJczXMlcuzHKnUes37LmS5kpzeEavfSsfsv2XMlzJa5ieMA3CLma5mv3TvJZPYpv2X7r9l+y2eybsv2X7L9lJpO2O8xN+y/Zfsv2WmOdYsH8kf2X7LifNmt7Iqdggy/suJLiSeLotYtOdc7WR8SXElw6s042E1glWbfldV1dOPs3qFqoFxiv+VxLn8o1KBpdrFVBLGxHo66OpBYkfSmFe141H9meL8NFTownLrYCoWRzfqmipgiRnpvBeUokIwzLovGylRFJ/CYa9jooPAjeNlOvAjek0V/OGmsDTMzrqylUFJetKC5nBRMGS6xTihNvUgvESK7dV5Rq0b+q/mSXgi6aMYr8KRxwXleS6SkoiHH6cspWRs/Ys167OoxjBcsnkzJ7cXTMUiiAcX5ZdmRLAxMx5mTVuyi0Bt2ZdootwIV5SnUACg/eK7xXeKLoDhLoWwhxEGPdl3ZOSLKeh5JDrReXeK8kV5YotoQYewXQQBhrQ8sV5YLyxVm+KtAYpXJeSK8kV5IryMr2j4lSrxqx8rLysvKy8rK6f7hZhKEI+Vl5WXkZOVlSJ7t/ysvKy8rLyqzZYQMP+Xm+ReVeVeVbpP6VifjyLyLyLyIs/V2fIu67rup/vGiV6R/IvI68jru6vVfbHRvyKu7ryOmJy3Z1YrEGSrejaj2dd3Xd1NvJHxnzlXvRswYjunnJd5I4Y2I+WzTQbDHh2kuZLtJGqMSXtWKqFY80e0l2kn5dnpSivbMBQN5Y8zXMlOHlb1zCXukEoG8kWnJfs6JX8q8NgS90g1A3kbma/ZTqNJ+tka9yUFAnkb9k8XknprraGvbeCgTyN+ykPuvT4XWzBexKKiTu37LiSsjb2OkWTkGuJzXptJRrjgvGyeEWTkGupJr1IumDCK8bJ4RZOcXPUpFGkPlhxZeNk8YsnsD58BioVEIn6surLqynaHGXiMdCrCAurLqy4ZFujjL1y2EIMAx4XC4RrsBy9OdlRhGDcLj6Wb8RzHRck/wCC3eYMq1LrP+C9d9dUqXrt/BpXHrwz6TUw/wAGvacFanWjUrfwbs+mdXh4g/wbv/rQv2F/BtDeVOuZrAP4NarIwadmNwD/AITPypDjN1fpyKqN2NwfP8Fun3lTvNY/hsUO069/92dfhcpnZ0akzyjfcMmfn+AlGLz9wlZQLAkeV2ZcsiUxSl7B6yDbFYbsy5Zcsp1BSl3OBBvBK/kZdouuWRKoZy5OFQ0hdmLF13iu0VOuGb/zhL7jGChZHNeSK8kFMFeb9SDXvONDugKvLFeSKIMJF0eK7GVv2JWvXdNGTL908pMntOu1ma8Dum7RXM1zNTt9X72yr05yURzg3BFwREM4kxbRX9Kc1GDjb91+6lN4M9whF6pzKApDbgi4Iv5iLdk0vWs2UMPhjxNfuv3Vi21ZeO5dYNX149SLqRcFRSOGHe3oKvTarHrNdZrrNcSRbRrBKmf6jdJrpNdJrpNXrUqypZ8gv1kusl1kuslZM1UOZVKefR10ddHXR08HQRvf1ejro66OujrotdnLaYa8a8a6LotsfOZRj2p+NeNeNeNEC0o4TdYeFeFeBeFk4GTi+16PSLrxMvGy8bLxxV2k4p1ZBth8EV68V4IL14K3lDsKtY/fxsvHFeNl0ZHpisxj2znHERY+CC9eC8EFOoIkXz51Hr2BHJ44LxQXjinHFEzR9mssBQGKcfDBeGC8MEfNAdeKzVQbYTP0ZdWXDIlcZm9UgVG4w1DpNurLqycUZM+YNnf2gId0U35+nCnTHJ2jYEmu9EMgytwy6otQRl6MhrvYEoXBzf6Wf/IlOMG9tnX86aatBfhcfQlgYl5DFTUnkoCgJvo8minutJRGcrDrDF/AayOu3nPYUKMXdm4+vPCJox7euWwhjgKP05R7I68PPYvKtSFW/g5VnQYcx0XJL68qZIjj3LrOEMK4/ryr9/1lRpeBcpnXK5TzTf8AzV1uGXZdlynktO96tTNrNTqdmXdl2Zd2UiMyiRj/ACDyRXlgvPBeaC8w1qmHLPy7Q3oeyJeyJe2Je0Je0FEsjp7sbgV7YF7gV7gV7gFoeteq5utAgHvAZmvV3Z79dk2hXde9XRbY86zHVqu33KsvuVVPqVWX3SorZ6NwdXZgGbbNN3+61F9zqp9Sqy+41ZNI46cwbdUom1qjv9zqr7nVUtinF7Vihbi2q9Mj7VSChuU5r7tVX3WsvvVN5OauN6+5CTl36YULdqFb7vXX3iuiauddk9yVZC2YTgX5DUDIezXLH7mJPpC4hepmlDXIOX3QaJ8mpClDYFNvusFZ068hivjJEGsbn7rwv+rKjEjqeSPvurVsI2BqmnEWoSUJajxaPyupIkdHu0zsZrBY1G+6LSp3/Y+3aLoGXqdHzr8VatmrvVDvWZfbr/FrPt9Y1NFkOho9JU7sGs6JhypVtuwvtt1W80kJNX1TvHMu8Eo2hRs6FjtSoa5W+2Wk+b6MoUtSxP7adketOvE1+3YJQzNDqbGlYhYCHNhVoaVgv2oiNVauMlu1dsVMi31lgRmS7KFJ6GZfLL7a6uQHRHC5f07dfKMwhYYwLSKKlLNyrPX7WyvDr54gzv6tyODAgGyRs2sYdSWdjliD7UNXxVs4NGN7Uswwa8X+zgWz4wTo4cRV3yK61B1c2vl1rGnaHh1Rt9orLbBH2A4wIC+01lvBr0aWFnvevfa6y+1VlsVvJqxyavD5NRfI6QK9P47nRt3Wx6a+z01ayBk3fs9NPj018lzggB8boBPZbJpr7TURModX5B9sqp82qvk+YMTfGAgkzZ1ZPm1UGnHK3vQrp6FdfJcuNUnxkwDCaoBEo15xrCjhaTVQJ6oV8ixPWl8f0Q24tXErOeCyGtJ8CzEY5NIEHbZ+PvSni7obaYUFezK98IiFw5jYRYFqjLDR+PGziZHycdhN1dXswGgNi28ZVrAbYz1h2R2Pj584md8jGWUeJNfyAX01m/kKpdBeHapBuDJ8fsZk6fyWLEHOJY3MUFyTFv5qqXgXY3M4F6E8C5myr/KZ1yVrobcT5dexLpeqIOmEkrWfXvRlgHpvHcs0Xq6Fa9EuVXJLpdrIeiKT2surejL46am/3nQzlT3Kd5SoAK7BsBXudEfPp6MX+OkrL39SgqvyGnZf2AI1YUbFrZp1F7964mw52HDTrUYPaaS8ZyqFMI3ua1Skvul28o/HyWnr069KEtAfPjtWECiAD29CvSi+5Z0HH8dLblXpgpwPoBFLrZsoFYNdWLgqsTfIS3SA+OEsyBWFWHb0QUm5vaKq0K9FEJAUL/ydu9f4/Y0J16oqg7NsNMfsXNZU8+vQbyMtb5OOsqWFZ1iVqoqopziOJdKxqzoZQM6Plh21t0Wc1KjZ+RWKtQVMK0dchj5eOPOjOyISv6oaNdvP8g0KNQNGvytrY9CGLkelGdgQ1PSrsO9dLq28imDPqstC7ChV+PU5TRLAwt9zrSfdv+3fwGBRosSMlKbRj8fj7dlyRgp6FeK+RXI2bHxiwGvThcDNd2dBk09mU4xU79eK+SWhHqfH7EK9xtCu6icc1vO0X8sesr9eK1ijvZ+Pc9W5DTBJo3gTW+CNqll6MLtKdwEFcsVbYI+bJt19gB4to13WoCvqU/j+v3jK2GCJfrTa/nEpHz/kYi1G0BqwSnfDS0XxbXug4lo1lqY/nNmbZKZK2uO0p3AEiQn2SVXaqWhy0qq18wGgqVnRwxt8iqzJ70VZAERKHyUBl91qLRHS1I5otWhOfyMAQVNaNwVqnWJMXyJ6ZYbNIiuzpXxiz71GxHTJXjX+Tgs2bNevaeWkfNYXyOgVrFmjbHZxvHLPs6gR6HywFNDvC1BOMtVC+Siio7NQ8bmfUtPnvsV5WNb1AUflIdNmC8F95LVkP5BSNO5VpXlWoadQwLFiMND5Z6V2ter3057YFL5CALWCVNCP2uotOlG2evjRovKzbG4Pu529MgI2d4bSq19k1wg/LH7FWiUrkrR9zVtS+z3TGuWgZYyX7uus2naDUsYtOw7UfFGdmz2jmaVwLUR5wdD5JVjLHo6r2nyq5IjyhAYrEqxri1rxKnx9qktKxTzYFNZ3yV82Um+01Wl6PVWbdohBfGzFJOo0I6m9UFLJxLh4tl1Yj+2hVtmpDDi29SAsqABaZqGWKB7evoZmIKnGVCu69GEUfz37dH48Kg0qAFvbIWfGyjakvSB1fNrrSgKlXycDs324CuvUza5rRtGzjZUc+q9EE1LOCzSoQ1NYeUCEfSrjXyvR4n8eo+1ouOM1KhXdb1cNXPzccUKrZ9eKk0AwKSR3xK/hzJVhTUsys6p0hE0I51aKiKEF8sj/AE+K8o6jxaSlRrzWtlhBTz6VadSIoQTrQrOC98Tt+xmyDCaJl1SqjTDV2/AITL5Fne5UzL75d4comhOmAi3MWAGznrWq3ClBpx3cX0SfGt7sukZqzk1LQ6sfsVqPHC08wWkJ2t/HLuPti1RSCIjXsJomoXx2mTty2v8AGIlfK+TGzyBMK0O7kVb4uD4yEWBoK9nh0B2Mi9hkyPl47C6CsRLhetMWl0J/dO3K0fjVe447mt8efN+Q09NrmPWvqQdDMVXSBc+lvPBejb+JlrzrfJ9DJnT26GuP7MOCd7FZCNA0XblX/jlO8my9fGep8y8cojzddpZ9qum0IQmztJiBgVrfxOqZ4R3cdB+XVioVOnab0LSteedhqLKxtUM9pa2joL/p72Xr1A1IuiXxwkIN28h5VWmr3yynVeRdjYVT4xUryjFotKTQb3JHceVI6IWtmhv/ADPvOOFobE6GPVzWRCwFGMrF5VsoIp3dCvnjt/KbOkSl8U7zEKAoqzdHXUc6zoKuANWGtv1syJbWj8nNlfH6+Y30PoymWlkxBPyR53Pkw6KpZdrfs0qAqAlKbQZym3SVagqIXPDt8h+Rud8LAe7MQ4igrNgdUOfUnqWfwylbCz7mpLYtfGMqLM302tD0q2RntnVHkzK3q1wD8krB/jtaFXP+mp/X67NwpTjBtrVDGgOHCqnDIf0yfza5UyRi3yC4E4KZGrnFdCX6W4eWthT/AKBENATfI5Dnaw7sczUHeCRc8r5JVlGNaxGzXRrAgtq5/BvjW2wBD0AEX4kxYP8AH78ZNJldetMNvKLCWJ8mhKsLTASNuoHRr1jlxTs/00407Aft9ukXL+UCsVgaoDDvZotFq2jMJufpr16N2FAOnlyp/J69itX1wWhzzWaVe+0yJ1r5ufbWZDWzXB8pryBDao6YI1ZBavoQLNS441M3PNLIsa9Rv+o68Bfcc7bYcrFdVtQNiSNARIaWNRlLHLsVIz+RjACvv5+m8bEood8RJ8q0KuYdvMqwlk3NYUbWrXetW+R0rEh6CHdER+VbHVKOzm1ml02UElsJrlR7ka+VKhP7mQan8howeXyIJCW9FhRL8ktWHw56Qq9rNa5GtjvnS9+wNF+RUwKXyKFic5eJtD5YUi+Pz1maeOKwwMn7e/t2hI3yCtWb761ucRSgtP5Z41hl1SShihdQzPVXnuhR/kA6jR2Z6c6tQtaGx8gFTWSTTuGq4FcDNmxCu90KsbnpwfUNskp1jAhsagM6NO3fuW83ADUj9uHBcXBKxsSpj9g/yAwg2ID0jAzxTu2LlzEwIUISzQuvXsiVvSs0hhKfftNC1NHrBEPS0Z27XxrJ8Ap0Azf1jCVq/bpjzi2NbS8Vsq+3CXyG41q98Wp+eySkEr+oQasWblUeGWxas+C0VNnBZ/lpGe1iQ8+uSqIy9F4KxO+CGPZsEXr2SKOcFn+RRjGjEjdHAM8fQaKNG9COVbsNb9Y5FCgGL61VrWeV+4Mow9PN+3wZW611xZNq4Cw1UhEOmETlFEwtWlKna+LabWq/oiV/Psnr1L12laaqQiHTCJO34+QYr1Z/Ht/01GnXmtHJLcrQs3syz6TlQqYgp4rb+PeRY+4XInSnS0xX8X3QWDaGOWFNrERVRhbhauCHRYZrvxuxnbNHba/h+4K6fSyD1wgujGGAm4V/Lr6ELWLcxpZfyWsRHyg6le/HWzC0vV0IjDAbcKxVFaha+LOCUd6zQQGo74r4NXLNn2KN54wjFkQUSxufFa5XkXTxUHTzdiFzP06sqpasnhGPHCeLOrvxyncRMjSzE2wAisjss9awESCQRYq1L+p5VjRBXc1q2YdxqTkazpaTUviEe4KYa0eeFyrV8FOE9W1fRMoRJG+S+OIPjuhqEo4tahH+y5UyRGx97zThhl0rVz5FSxw9dP5AfL+MgpJotH6OrOo0Z1Pj5totu5Rwa+p8lu7Rcn4r1UBtBvpo64qSpYtjcLGIqIN75gsvGsaxKVEVIP0u3hUQ1M8/yIgxxAPa3BZQTWLOxcw8KGbDjj6Tm0Ilcnyi7XrwqhnLhfJt33CfHMf3Cs30k63jz0LVCnGjWdfINL7fRG3aWRR9Cj9Pkh3HQw6TUc9Sdapfc2/iYe1pvpcfrV+NgYUPp8jh3zmE3hqS71vow2p/Ifo606rVr3wy7wRlwvklOVS1VPGyD6fIM73KoDko2c2/C/VXyHG+4Aw9P3Q/Qo4lht5Es0/xr5B67xlytHNFpV6tk2RYZ/o7LawI3mqWrWNaxt4OpA4h2oGq2vjtindFdEuFaqDtC0/jZqT4ny0lVDNX0q9nEnTsVdjkv04Wn8cr6CZtL42bN+U1tKN7EDzG7az2r2hWofSzTFaHa+LSBIXyG1VVYdHbAaV/Aaju1rv1eLOr3xyndT0dTGfP3ByQq0JMTW9IorA7EfoemG1Gx8Vgy8uhktXNSuy8ZFt/JQU7dPTfTcTMKNwd2wbMw6I26tFdk7q7rV6MND5UYqyrFDxHld0RRxOD59SoEX9lyiFiKOh8nEF7mhYtzDv1RU3ztG5Xz8qrnyC4pw5+lvRDUR7E7SnsirzufLp2mN8bsWo586uZCE4TjypkiOJNI+nKpCrXj/1i1azd07nyOzD4uwULQGJRm025WnqizRVMuV6ctPkb/MZhLXr2N25TynySC1Rc8s7PLhaFwu7crQq49exbP4bXyUxamLkvpGAE9AYtAUpdvxraEc+p8ZznEMmhBn07FgNLS0i6csDK9snktV0K+Iz8q3/8hvynEUHvuVbZrFKnXd5S+O0ieBrFgCDcFYWpLrn4jcQNbFXXms2Vv15AHGH6fHGLZzvZMBBsjO2//JO0+Yl0Rxl1t2V8ioNUnA08+3iPO1ntcIFWIC0qnx2y9csiRHF9DyL1TWF8hyo1pVdItQedOdir7viW3SelYpXIXa5rIq7PbOdfb2KtrIfPIDcNFUykMC/614Ve2XGsNLlj6IQu5LdpPlAm1/MPjmb5CcljP0yWwWKjRs0NaNmXZmYmoPnpbsqeLVmEte/8flT2iQM3GhVhaPlPTvhvDLZHXi+iQ69GdhWcatZHcFqZlensFqkFOFlVfkPjkM8CxPoArqVu1aUcuMpWMkB1rUtOMGPxKjs2qkaHyGtcXliyNrhjKXuXEDMCB50YOtfL0JOO6agWl8oJGNTVr3GnZENT2PIpVbFxApDrR6K38VPc2M/Aq0HYbKUWRc0fZ7d2mzfL60lpfIzlbuW0Sl8RMd6GPWoLopMi5w3ka3coD/6u88LfkIiXVn/FjW3oZQKMeilFkTNh2t6drKH98ua7NTDmwv7UjrM+NEtvToCpj6qcGk086MHvbdjJUGvb5iirUA6u9O6snEJoSp0RUxcKcGk0qDDe78gsZ5s3JtmNKgAS3fkktBZucTRNTpjph6og4kZ6bge7sXLZcnFPVEMAasfke77pKdSd6xTpwpgiyMKJWnVnXYb2fkV+Gf3i0Iij8s0vPYhHl8qn6NLhGrjO1wZqQPjwrFt4Z8Of7L5pYX+mvhj8efwj0xHWyE1WrlCLbiCkKv8AT5P+KozRhP4cTmoj0RGfcrzrjya8rtIYYBityv7ObOXcXw690MyNniI+/VLlWatQR4NHj6W60bde2CVQ/wAc2vt9hnaTXcmBhFGbCv1qgYLhOjBicermzzT4+4TLLKYtilo4IroatqdW5XrjFHhcIg2JHZwXqKjpEzy5+rX1g63x/wAyzbkXsChGMfpKHLavxqJVXvWMg9HZq7ENfFJmtjaNfyR4dvo7LR+PAuq1TtYxq+yC81yiWs+Pp1WeLM7fR4q9jV7qv/H7Wc47rGlMZxFy9moRo8O30eKtUA243fikoOzWAEDKQD5+7WMoSabfS1Bmtdk8lKTRa3vBEr+ge49cfaVL4bMsqWYGkNocLlPJPJmbQ+SAryukuaSawOiSp8fuak8zBr0GYfC/snknlwtL5EMDxxjXXHsxyaMQXdqxk/Gw0lGC/sndO60t794fHpTlo7AMkN24fRNjfGXmhiaEeE6da+08J5mCwrliyOoLb3CaJMvNJpmpUx0w8fR1vazhXxnG9WfHVvlW9woczlh5bZ9eEU6dfJdDwh+P5jZ1B1r32z6cyOWfxyh7Fxvo6+TG/pcar6tFTdfJLHs6/jZy1R+OunXyH81MWHSl9PknEqzR5N8Qn4yN9NgXep8cl/SfSTM6MDw2qdiVO4E8CRWxRa9S+MWn8f0dfKKUZid3Z/iux7IYEiRfJ82NylgaEhE+jsrlSFwGhSnRs42tPOMG6IgdTNDpGzdIuWdn5b6PFbfx3lAIWmbG3x3YX86saYrNr48SvYhZH9HblaWSHRhex7GWWpvS8Bs2tsVx37WAelohvj+pQsWOh8TgRV/bpTHdpa8YQu5Ko7IL305+jw5V7DrXlcwLWbKM4GhUsWKirfIhTYZolhz9HiiAgWNv40Gas556r1bB6z1fkX4+5BVyX9Vb0gU4v8x/nHIe5GOMckKlAbWK1QQB9OFzwnkpS4Wj8gDTY+ubUmCPCn8dsHhjU6VMkRr+yeS5V/VBQjobNrRWfp0KIZ2Lu8V/ivhjmnq8NHhO6d1atipiu6ptRCuwzHtfJu8KOYfXLXx/tJqdsNtk7p3Wnsztmo1Q5Df9Qepe1tgmkXHwnvKtGeTCucViDp3W3rtniyM30x19J4Cf5USA5u85YuF/JjdJWeBIzg6t2YVQZNOezes3A0o6Vo/p6WuTSGKH5z8qdSoPQ8UueU6J/wDJb7N0iXQ5nvELQrj7WrcGnKwKkarAGhGUlu/s+W3WkU8AQ9ixdW7U9UzNHz1n6aviPTavdHYVmHkr40/HoqzfHXXhsXVv02oaFmDRJ8csexd8limgnHYhrDfG2oTacZSaLTvzsOLOi8tnP9G2E068/j9p7Dmv8i2c/wBsGJqtoV1YtDrRkSzeT5gPBo5886w1o0YYx2tSviFpQztEuVYjLsys6YwS9Y917eOC0C1TPmWCaVmcs697YepMoudqC0RKUmgxdOR3Fndp6WIG802uY5PuZZIBG8ub8jabxm0mVq8KpGfs6KBUhXhfww21cFoUGewSKzfkJINU0Q2/rb1RV5PXs30IEBDs4oyrUz7USV9O3kkofJA2WGWJGUpNFj6vllDNkabii8CZA+PsxV8k+TTHoCDc2SZ/xSEFXpBrLojVYGh6tjOevsiNLuztc2Q11p/JJ2FXqmvkzvivDV6gq0eisVBng0LWcga4LCPaFXHc+Rzsue03LBkaeZ8YeSCCAYdVaoisxYlvOQNSvabV3g57dbOrOzoMyYSyfj0joYmHHqrWeM7tds0VDUqlhrbhNEmflPVr7Go3DR4WLhvbeEOG6qxnxlNtAtVX9sFarlDlasxpOR/kGk0ycLByfdNGK6cotBxz+7eBbuhHQsUHLGGXnxi/y3T9g6+P0vausykNptKoSo5tuAB4VkdRCEXRgw4Ah8xs97VPrB8ODGMyNXgeDjsUVf0IXbVK/ItYWd+/C+S/gnlaNosuuhFWKY7LELZoRa8OvfYlq+q1IdZuF8lr+fPlNzBqGevYrmjYDbo9m17E7dDG2JRrtTJbeI2gzstqj7tR2dnrHnVP747lOdKQFbkTL0g65dGNehGEuqeKv0YXwWqpKZhEmAmZoi1K+ljuUGZuEzE07Wk1amOtHhPFW6Y7otLJJnEHKQZ0dMOlC7n2M0wflMyRjVLeQxNBuF1VisOyPT+OzrKQeU1lpNT0bOYg7xtGdbOjCTRXVdVMbTjf+Nwm9mgSuQOg451/kJhAq37OxGrRHWi0V1TwUo8tbwgmjfxj58qO2atL/qQshhCbTQa8RR4XVdVwjfEmJrhrQCmgmZf2TyUlrHqygOxKuxymtmx/jEnjVpjrRaCZvpJ0R2Zt3VrFfwuKse3M7ZWWW8qGSGg0YJop/wAKTo04jjt6Qrh6cAgFd1iXZ14TsTycCFRNFcfR3Vs464rp/uNnNo18ypsfIJWpLDwntPGHDM30ktO6OjXo15ad8IIVh72z6sOXd8+jPQs1q0KwosnTr5FdjUqfGaDTnx1bQuPkYsiyJKKwKPp0Wb6SXyknKyaPamzdWmtaz7WjF5Rr/FhT8rfR1vNJ9DOh0op18pd2U+72LXaJgS7DTsturKldH+Yp1YD5wRC8CO3C+I3vLWZHBGKDP7Zqw/t9OF8izPXPwse61c8Z9m3azHz82xPGvwfllwnZa+VHRCULinXtTqGytOGgH5Bm+5Yx9OeaaEmk30dkcEDj18KVF3/D4+67K1jl64/yB4PGTSb6OyeK1Pj4rquUi1C51j1iSq8ky/kTO8ZNJvpwnirVQdoeh8WmNBf1kI/iJS3ujDJAsV/dOyeClDs134vXsvdzLFFquoSrKpvQIhlgVvpwytQ/q+vCf8KU2Zcq1pirNo7s5KZXIs7AOV6eUCizCTR+jyUyNFtHar50bd23rJphqRgxrks34pASGLqzR+junkr+iKhCzaub5JxrZUbJZ2yZ+KbRJnZYs4bR+jundXbw6IS2S/ILpKAaedp6k7UfG6wcDzqMeEzfR3VmzCqGbm+RaHUFY2xpRoANKZiDHKb4+bCjUhFf2TopGHAbS39WlDpdaQxz+T6XvXWWeOE7cOJMnUlz9y2cZv6GT8Nb1w+s37SM/wDKxbwa84/XVlzogbgKJNhx3NEVyZJN59KTOsvWCQKdfJYctkF8+d9LFkdWO5GAdWzHieBd9HRqa4LBrMeq0KfmzPj1726P0daxI2R2QSATqvj+rEta3pQNX2strtf43qdmb6cKTLYpQ1jzDIc6VolE33QRpWoi1o4+vOgSL8t9HZFjHrZxo3bEwSFLM1yVH1K9KxDN1z5cq9kdkf04TxWgCsQDYM7EW8tMkZj0I19MuMWjpCuwZ+fq8U8VsApyCHFsuLrOvKtZJWNP5U7Qp6Ibsfo7LoniztsVKoUHCM1dp2c5627xA/yVol/6grK3+LLzVzWDVbT3p31W3LFpmAUsqeDEbnzZVT0NEd1NH6PJPLlXNINOOxuz0JUJdmYhbp8747ET2c6Qy0NKFmXVcp5KUlo7kRtaveYgtMrVghlbNlfH4VFYoSESjowtfR3TutPVFmjNMmoT7jCqi3z2QwH5JY2HGjGdIlSdK+O2v7J3RJxHDQuk3blUbVq9u+/kMUh105fDymoV5Vi05U7w7UZP9Pkt95Pl0Wo1Z6BIl3DeKMuZyHHhfHKHip+uXPerbHbg61bXqUcGt4qtc4s/Mix9gnyg7yv1IPIj8zv4tWMxeM2Yq9kdkauz5uw/02rg6kY1CXpfII9NexN3JoS7i+HRganwbNQjwsQ32/qvjRP6NWb3Wdeh1lp0I1JTfy118deNum2nOpKo0T0ac/tG0yd2ixLRb8q1SFSHyXO7xX/1k3G7RISgtqj455GnHSqopYAg8jaziBAA93G9uPClHs1a9IT3azHBi7MqU2kzsrVsdQfiNqvAURR1ccehGxUnVLIfZRsygqlkubLP1B34c/S9ojpsOmS4Ro9VfzA3438gufP9LDN582WZ8gidhkYkfpd0/HKtnu82jwrNENyNnINRaefE6Yx84+b8h7sGxA7J3/FzTeRKeewpdUQUSI2RGb2MYgo+qda+mKrZv7syq1enalQxekq2TKKDWGBuqeCuZsLCr65Kc/I02MeAI6XyFosQ59M4KkKbVMazoPXqCqw4XVXc+FpgapKM/I02s2x1oauy8okMbSnGDAahmH0J0M4WeNorpyrmfCywdOdSbTaTa21CkxX7OUs702i0EOEzExsZqMGiuqu50bCDpzrz7t13Nj3yY2W8gbunF03Vl+q+OZPZ2ZdVboMSQdRxz0L8KVTJaMjNE+mi+KnUtWPaP+FnU/etRi0W4Vqh3kDS/f5Ib2CPYjVrEqSmDlhVNAvnu0Rqi3exkD6UeOVZoO0wabSnZftM+zFpVM9gu6+Qs/3K52ZXITcHwuXBuFoRJV0Ld+N98Q8a117JdGVWpCrB1vVpSLW7QecZNLCtPU0RfzLJahKstd4Xh5uuOeawi6bwG0IuyINiw06cqVv8r8rD0fbBYqSqsC59svk2a0BiqFuzjH8cJ4rfxufo7LL0Xoy08vgeJueqjbQ+1ahKZGjwuFwr+cLQHezyZ5f1dQLKnIU2ksz5AMkT6/mlToMJ2guE8VMbTjpfGlGfhkWHgfM3ZDlDaB4ZaJ9N6dGFaDRXC4XVXMivcV3MnWgSD1CUNWUHqbrTgS0fWlUpwrwaC4XC6owImh9trr5CZg6MplvlyfjDCjXrwrw6porhcKSt14FHAxM4ulpEmzkeyXPzZW45+FXpLhNFcfSatV4mhKwejc0dOTLt7BmlBo5Xx97KEGAINFcfSatBgWB9B6Fuw7U2cvtG8kUKErBMnIhnwZlx9JK3AZRWdCUTYmMx1ubUa8fJyu6xs59GxGDRZmXCkrwRECSx5jZOVAcf7N8j0uX7KLr4vS8VaKZSV+uIwM6XltUqUK0YQaZN+41HN5QjtGGcZoRBDxhTstuhG0EBfJWpZ4oRTr5aRhWzWmMp3IzH8SN01oq5XaJ9WjA4s+s2rbGNoMnW8Ltn+RntFdu3ZmWZb9ymtasNh5TtU1of2+jst/O9yq/6v2Va5OoelbhcB8hoCE+DchWvQ/t9XZb2O9WXLp5SWTsSqk1xBAbC1WpnFJpRdvwPtxwuFZrDtD1co+bNykZQnMZBjnfqZGq+cQMokg304XH00MoV+OhTt50uH5H5AhzL7CgAsDQ4XC4XC4Tx5WniNahYz7FI3712q3XgqmrAijKMm4XC4+nC0vjcr2hSyq+fFoLquPq7q3pDrq3oEsKZCO9yHtvl/EkEURQ6porj6PJGNEI9DTnbaHZ4aHjNINQhiY/x2FNcJmXH0d1OTRbZ3J3CUaEaS05RsG68PVrztlycceaNmTN9HdSdfI9rvLKy5XTzt/ZKE38hGaKqVHuno0h0a7N9ZL5To9IUsmRFlk8lLVvNRqzJ5Z/qqNT3LIxMOEW+jr5LZ9bOqUpDz682KEH/AJHzW0m45K8Y1sgXZN9HWm/WmH+RXqfmadfJndr13s44yn6+LNx67K7/AH1J+Otny9K+30dEh5IawSInYwH5Xxi3wVnWp/NfVp9Y5Fz3aP1db+c9Sz+yk7rB0XpWLEfcv6+V6xfjmr7Qm+rspwaUdvIlnkk/K6LKvxg2ljPXWFtSpyjLllZIQUI/s3CKJiw2sGVRdFWP4lOI9AVK5Zwy1Lwrgm+nC4TxRgQOPT+LuJRl4kP8vR0n8tPUhZbsyjJpsnZcJ4oteB4X/jbRXiIMozs862gSvKrqjM3PLd4PPj6XP/K6rhcLlX94FA09IEVb1yWE/wCJE7PMWY8rdDKr58eqaK4XC5WhoQphD8iHOvcszsI5hs5SQK46EpjzMutQG0VwuPo8kUsRx29yVlqsatIFq4x3/VCrytE+OAAALMuPo6dfINv1mCD81tekCtYsSslf8r+yxWfLjH8pm+jrQtxpVgPO7aC0aNSnqCrT3rz27P5ZQ5Xx4pPNTtQuDZcJ1vke3rAjzCqaNFV9p2PsaH3S2GE5SttN3FeehYqXCQKyduF8nM8aQIeRsab8P+Fd1ZGtaunDRvWxz8IgykDu9OzW+QkOxCwtVz/1F3SG7Hzz+zVTq7bnImjRkM9Zu0CD4eoV6tkG2K+9OcgW9APaHxyz6V/6Or1xwrYpPUzXizt1XVkP5BOtWDZa0Iwi5d3M0IaNb6v+FaI+zLVyJZhuGX4VTaerW7wvrE3PUeLs64TNwpn8ZFfuSKS38ZhMBReEgjeGQ7gbAR3Hi+RuQtDb8suFwnZX78KIwY/trRwzZ7wt92gdmY29OvLO1JZhKl4duK4XC4Vk8Kwx15bNizkdoHC9BD56F1bNSv8Ac5SsZ+/E8fdArTf1XC/srFodeOx8jd4xsyiSjnzDCVuv0r0rOqqWTXoq9RhdFSvkolZlwv7J3WjrwrR0NKV2VelIkzXB1k5XLLKwJcuCDw6kw5gLA4/o7qwaII7u45XqZ7cWLpSrs6rBLbNm5kaAr2f5nz9L2HTp3W7r+iMcZkJcl40MPRcSTtJYOU9w8wxJCJJ484SacXTuvkV579ymEdcdjnoXyWTdHXR1P9I/G8/08+zSnEtK5G5BHJEY83mxY7RAFgvqG+RfkvRU6/d/H5LwakZ2bFWFsVezOqTlbkvPKvD+oq/ydPY1iHWeIUhVxR8xxQYAIQcVobRJhn8GaD2MuFCTFr6w+VjF4mtC9Jp0aUaY/kddvJJmDbsjjGX4Uos6zHjp51c0oy1AyrFz7cb1RX7vrNRo+BGFEsL9J865+GXLLlljWR83a7+POvSxrwiRLBSk0WIYmyQNeFcdupC4C/TJn2OzLlOzM8Ce/DF3fWeMuWTty127MxaVKFUbstPLjoQtgJTNA8hSk4dJOU1Q2Ru92EVix+mjoQojpUZzKzcLjlanx5rD+WzRnGQDiuUiVGz9GUXobXdReM24VqxCoIYybJhwaLcKY2m1rGecp/tO7ncPXtSAT3WTaArduUoxa9uxEr16TqUiXTUa1bJZrE7FijiSjKMWi3Cdlcojtjp3yZZmmzsUzBjpbfKvXXNPLpwC5tCbNXCW2XLxo0W+jx7MQJMglW4O2KTq1ahXjs7MivQp8I9ghn/Kq1SWzZ2dDPFwnZXqEbMaGpLyO/K1tL0ASedqwb+gHEXC8brxuqOfK9ZrV4Vg8Ig2m3M8WcDRND5BpejUqQiCNCm8237bmJ414kwlk0vuOk0eF1Vyk8pU9BrTfKLfhz6I41Ko4y1SccNpk9i90VUDdaI/JYyQtLQZbw52Y09idFaDO2bWb+quWHvFBXiAdCp4oD48pHbwAdvHd47fGXZ1xyxhkoFOWFyrkdpA1tf1lh1fEbha4fNQ0XZ0QncHZdl8fueK3aqxtiNJzN8Yu+Cxf0IUBUKcoy4Tr5Hm+7TafaPkXkXk/OVcHp09OtOoX45reKcyRHGZCbZAhiKHCdlo58dAFkM6hu67KX6yGR78Mbcau7Sbi7oTsFpUoVRdVwnir1CF4WjnlzitN4vIkLsP5lMmXtOFVbcLMdPVhSjQpTkSMVwuPpdoCvCv5FjLkKyMit0515U7nZUNSdd32AtXCMuwcY2i3C4+jxVitE8D5PpK9RmdurrcF4Nm3omtIxWC1mxK0SiOvUDVzbl2IKw68eFx9OFKKv1YWhUrtjNle0iWnuW+Vn1Bo1uZVmZJdKVSlCkLhcJmXCJH8X6ZaRK+8xKmnqOZVA+yYj9k8VUozuHz84eeFm+nCky0aULYx7NnOldMS8dnjli8UpP4XXhdNXlJ8bMjnV2+pINJrcTY09C3PStY+e9sunb9WtKMpy8S8SL/ACo/FM/16kWTMnZbApeY9o2ter99O5GPEbpvBX68rqnbx1MuPI8CHNqK0VcrROMhLAi2SlJcp1Y1xuqhm9eEuDPP+TSNwO7Ps/xqf9bBTblr9UleQ9YlGdGr0VP9TupR7R0f0VUn6yk3PdRN451LEbVfapewFzlEqMCXJ1JdhJ2Tst+g+bflPh/Iy7sql307EmDsUi1TVTUbM9o4BNCP1da+W2iAnYJPIu7KU/EQM/uLT1CijlVhhAzcfwOjgjYHq5JM5+6tGiYYiuJ6V6YXzK45HjDj+DhcJ27LT+ORK8puJO/BKh3lEc/xSv8AVCnEkVwuPq8VezoW19ggtSHbTLKMFpkgRY2fatWaGd67fXhcfQj9I6GvFTk5HtvwNAtF8eTglMoxaDJv4Jq/dgKJ+1trnPnrTlBd3VCkXQPRowoAZv4HV2xGsLQ0J37VZ2r1DnJaPGMl43XidfGcjom/gkvlmh1ap+jUCjejt3Xu2vE68LqNaTqrUe/eEJgjZkyf8NdmzNUl2niEZl/ZvkZetLxuh15EezUesOrlkmH4tUevXitB+SE/toSjavhn6miP+0mVaDeGIfMV85+gq/dz1+iwZ+PUj9NU/ETBlXVE7HHB+sov2ivklLjSg3iskh0f6fGbiu3YijZrSEXB0IwhTnxL6Oy185tGnxKK7p5qUlhanqH2B2CTAedU+ZeHfq/w7uR7w3l1d5sifl8+UYWtCqDSWHsyzDBJEkHbhf3+rqcGJHZwZVUXq7cIfrwr1bLxWbrRJFv2bjj6cfR2+mjlh0R6eIbOlRcMWjYeE4E5Va7IE6mlGx9ePq7crotq7FtYAZtYB8eJbmKvAMGj9OFx9bV4dWNzTJad26xlYBaibRn4w1JWzYmA2ezLquP4O3C0tWIVZO4ySsgrIzxLOLtB8uiTTNTpwpBZk38BiNCO3qvq2MzJacNS214vRmUeF+ixcttCxGPCZv4NC3GlWk871jKzGq1Lz/a63X8tBMJTaIh/D8/hmZMy4VsrDFu3J2A1KfEbNPytUu+RfI5+S741VrSnK6L+YOjLphC8Wa0Vb/JrliRZtWaF0IGlIJJUJO/LAjKOeEMnL6hHHXFKT265Gjncjvwf827fRxVPE1wHaoMbyFVssdUJ9oOvkoO9fRCQRJRlMbwknaSq2JVbQACaW3U81ZpMK0KZKT07MLYeFwnZfKc71zP2dnlJEk7rjlYt6NwFrKlQs4+jLKtwnGcf4fkGPIjTnJcJvwqWoZ2u1RXGxNqecSBIzjx9OFwnZOy3Pjryfjqg2p13jOFl4Facs7Ycc4TgSPP8DsuqmNptp/GXd5lKNwlCFgy8sBkeL0dVxoJo2IvwyjJps7fU1EmpsU8uvRXC4XH10dAedXqaIbgNDYYCISdmcWizmIWuQhTmepRsWbNLPFSHwosuFx9JP1Q96oed7Sd00mmp2iVWkUk3d5KNKxYhk+v6PCZlwv7fSUmW7rPbfJzfKtTTGWXkinnF13ZVhktkwiQlR4/gKRhQ3dZ9OxWZxFFcYwtS7C5afomeKH45OZ/IbHsyqtFkzJ/1a+d9Emhxa0aUOxdK56o3KOZbpWsXGaKqDAidJ3H9YcJ60q9CnZhaDqWZEtDBEED920KHLieDTiay+VGrszrZoxQcrBB1GOMnsAh1G3Qsb0bFjNfw2HZWYvzkPzULX7vj3O5zkiGFnYJpIwYHrV2Yg5B4UoLoqu56dKtocK3T6yxrDnqtGdYlLTHbXCsmhWE9A2lTH+ryHJl45LxSQZFrlnq1z1rQn7fGtOcP4tW9IS1/jsqYowmuk08ZqhfNFavQAsvZLXPCbEh9eE7LTvRzwf8AT87Nc9Y9ef8AMi4bJyt4vC1fUJQBZ1ibNDI3IWR/3/gdlKbDjAP363ofHrAJNaO67jaHDxQLsgPV3vuw8rXNmEqXxXIrhbEJ4+xXPCyJcfXS2x1WMYuzbsaBdA/SUpGEYULJfM8KkyyzfjgAR1M32oZWh7w2ZcJk6ISMI7vyDiIYFvEhTnEVo5ZLoReMizswt89ekOqCXOFdj+zfR/wndbmr4hOTwNTJbZ+h11OniddDyfAyfSBpVp1zVLQ7gOPpJ+jbmo8wi5HEbjzqzHNbsckT90zT5lOYQfH8737t6hG7Xyr7nX9lduS0JleIoZ3JJweNGkIbzYpXun7IX5cJOkKcmeybwnhVqQq58Lp8aYRRFCf9uO9+k3AZSaERM+na+QDg4wOGKiUHWExs5p1njNxqof1Ld+o5Gp2mtgPH+bm8DsIgu6t6R9d64YSRoVASDKMDzYCl41+idhusyH3KgX+sr1Cxp32/LNCPkaTSga9DX1OvDfK8v1bDsOceo11EuokSEXane5YwvCXD2GvD+ujejQr5VCcFKDSbdw40J9YJ4RXSKr+vOMwEpTwNtuIk7sv7rhWrEKoaIZ6dqMVpZAdKF3OekboyqkEJ+pLitAlQPC3GJc3Y4aE4zjwuFJ+GuHfYtVgRCPhafx+vdRapM8gjnOiC6K7S7Iln7iOjb5ajsr3grSG07AbD/H7kJtOPCMcYIaW5Iqv2usYTkeNamOgCWlQKAlmu6zsttSedmDzh8J2WpUIIuZfHo1+Poc7VobGu53fvo2q/r5LWT0pS/pl/TLKyB6hKtWFQKsgjYFmHnm2mX91J3itTRhXGbQ8lgMHMToFdBLxiXQS+N4oyyd07fg7TxbY5sSCvO3h0bHvWqY4lIWRL9hoOujro6gGStP5CfGKHrVP7LQ8j26WoPSz+sYNuWHHTpgaAIt92tbknHQ6EXQqqhsKz54Vsgdl49L3Njlns14mHm2pAJJD/APKrNwG6V7pxiYQ9pp+EPuKHv8cWInn7zxsxsdn8qg/eFqL51krtIYpPHTZadt4qnVasIT9SasbULOkMwzQnYIIvm5/mJ/Isay9a7phcL2Y+QebY9qqtXXmKvRrtWHVL7AL1ON2tMZM23JpsuZp3kneSJDsqZfuFeoeYD07Q7gGRzQrjohnqWmjx9CiiWGvlEzjcsndl2aLwIO6Pl6ljE2uYxePDKTtFiSlvXBD6RTq5ThcDp5M82XaCBb6O1ilAN2t4nz7aoaUq8q1mNqL/AIWxoTMTOowphj9bNUdoej8dnSatYqxm96vZLq0XE9U/hmEvePd1db+qu0YWg41+efYuaw6sbl8lyZysGBSOaeJleITyv05EJoGllZNss4BiKLN9ZQVsc8i3WswsiuWx1h39GdqV+z2fHy5xpntaHH9Wv6pZuddulCGIYcLhOy1M+N6vkajmZ3Z1oXPWHr6L2J1QNYJ+zR/K/P0x8wmhYaLDhwnZFHGUKOn9puOVunyLRZmrh85dY7CFFgxbkS5EmcK5GMWPT+4XhDYcLxPFWlBFlPNsDswsh0uLWmYs7NuvXhVB8jsCkbmuuayA9FXJ1WDT+3sMDZpTWP8AP15bSp+WFC/7YavHN2761fOpesOTfje8fhG1NQagn9ft1p8HjXTsJZ0u9Ao2LAM3plO7RNeuxpgzq0kzfTcEE9S3ALjqOKQywGuIriK/Cy7Xu0tCt9ruZZmrW712NStRFKcoMsk3UrwZl8wyfMIMokg8V1TxTxdfzAkP0uBxNNwGcjNC5pPrXa/Vx/ThWqo7gdKgXPscETxIuCMjwLpCrnlWLi7DJ5cx1NCWgalVjXCzLj6OyMCB4bGManPqZlXsWa7la1rhsAJRsUrXkhVtzBK/tTankUPXhFlx9eE7crUxI2ovLRzpBhZtPpU/TsUbXVeZW2/qjyiOOmUVgk5ORyT6NcseWeQwI2LJ82cghqWS53xmtUnx9GXC4/LsjQ7xH5ca3buTtzv2vHHPHCdg0qEn/pF/SLJxwac61aFUXH14VojBHrMTz5nyNrYNfS8jtGdgg4NAfVcLhV68rB8+iPOr/ThaJf1v1mMOhvFpxsHJbsAi2fUix+385cHXFhQFakrRpGl8ToOIEWWoTsXr+LAuYxtkxzhsyaXx+n4wSV0pzW/6llH2kD7gy0TWC2KxNKAs+ehO2/7TZEh2bSHOkeseX23KFKzOP4Z1tsTxDe5xCV9Fez7be51swsupMVYknlmstqr5azHIbKqeTSsjj1b6N5JwII84ilOvZMEqlCXPEl+y+OW/FY0qnuU3GcBPMTUtQr9hs3DRfpKuZrISjYkNijPH0Gi849V1TxZSgypW/Qs2K8xmtaJZipVmCPOP43+rstCjC/Xu0Xzz8CXAU3ii9xhdqVqQZz07JaGE3qtXmxY8fR/o7J48tsfGojT+uyjIEVdlVmEJXFOubswycKndZQ/LLhcfThcK7QFeFp/HWz2NKg9Zvw/sOtfRHVs2r5LUuqmr8v5ao6tmFWiLRvzq1IVocfVlx9HWlpRCxSysSPPox5PIufcNXXtXHXnurIo3bxRiiOP8BJsOJzeV77cIsPTDcf8AmAJIRY2DSXkKvIVcld/j+XKmD+64XCOXwjnzJ7M4dLNjz26TQuravewaMuVyy5ZcxUJ8NSA921UB64JSYcJS8k0d2hHasDJOFhwU8vYGWOpaiCj/ACl/JTMFOwWYrR79QM3xqI/cZMiliOOzoMQYpGhmZmjEUBHgZnXyXp4WiB10AoRHx46/DxCyfwr4wSMq5rYq7XdWZhg8lgORakFhaIZppM/0d+ktCjAF14uIjiG6eEGX6L9FAvhKfXnGrZOWMq05V7grs4tC4GaZ2dZdrxFdfJsltGlX6p4cL8KfKdiJ/wC+IR7TaNedc+RqxmKCpWfI3H1da2WPSAYJgF/mKTT4Jz2qwlM8axs6VYn5qXGeQ5sSP04+nC4W1heWMo2IvYaa4QqNoYa5+8YOqWhISAWBo/wuyk3LbXxuNqNioWqTha3M9PjhS/DFuQmW81Fx9IrG+MPYGAMQDZv4OEyk/VtPYT8klYI1eA7dMtcjC7g8HLeisfBr6iCGABfwHuBrta1JWJHMWQ2hCqwrMQzvzAQ8eGeEwpp115K6+N5IbUnXH0/sr9+HadgpluHdoRh1iOD5OZx+Rz4TTXdCmtI8Zy+G0md4stQvUZLYwp7ByqVLlHj7V8Nf2tI+cErbUnq12kVdjoMrXLmtwhSY3teW+qhTRqvowX9UZNnwWyDrUmKQ8bNrM9KWZDntcrLYIcgAvpMzS1FL2vbg2r1sPo8T9pfHnK5xZoou4W65Y+l7OC4r060Jp6HjUS2gqWjDraPcMPVhdnDMsWull76l7KfzonlXx0/nr61Jp05jlKOeT26068JL0Wi7e0JVvknSP+uPyjJfPuNOxYi8LCeBkRiMujuqLlCa5n+3S6TqnrjY0IXTVpUdMN2H14W5kPoBmI8JEjNPH8ji8Z+MujXDYevIcWOStOxWQdkE3Z+y4XC4+jstrEbRa1WJXNEUVWJyvCGtGubywi/Kr2pglVvxsMuPpx9HZOyvZIdIX/R41qt/8nEPKuFLE8rfLt5bMsr44Ku0Rrj+F36tY1wjV7WIduOX6oZbdeRrVsyl7C/nM+HnHvzGKIofW/d9RinuWVCoPl2cKsW5BadQtpzWNIUCCsyXjPyJrajC+s2leuWxjiAf0tateqrF+1dYdaA3sy9QU3Lcs5lBrx9Ih7ViQZqMSMosdRHZX9VWgABLtjMqepUv68qhjezeIOrASf8AVaBfBVyQ9Y4FWLzItgrn0WHNMGaDVm6sBIEGdWkRNVmhVeM4YoxXCduVt8OC0HtQox4qMpr5DCDjFWr8etVXiFGwOvU6mrU2aQwrCcY9Rv7u34nGItQsYh2f7rhcJ4M6t1gGoGFmOOn4+5RUWUo1l/IUvGsu1Cldss3SzU8M8gsK1rldVwuqyz+UOpnx0akw+pZJClCT+qpeJN403gWVcz6s9GuG+HPuAoEjOLsSpEiFcuUlVP7IH+jr5D8fhbU2Cz/yl/IUJ1mdj53WodyTpnH1bwkHGBgvQukNJ/px9JMtTGDpxu0/t53kFCMGDw0a8YC/nDaShN4PS0p924k304XC4XX6XBx+6XB34mK2iVVMXRtSo0IUxND+DhTk0G7MzX7AywsWOXaC7dCWa5oEcB5JqZF6RHWP8cLaIMcRwZcfQ52DGbuRyGiFptDoWTuo2PIrUa8H8YXXhAnCBDDXUK1eb4+bDMq8crhXC+IQ64wrhdoutu2M5I051VoSq0q3SoulVPCuowqKA6Cu+IC+N1q0HCWBAkn5jM30l+i+QGE6YHSln3BADasRCGUwSkz1V2p8DJlq3Kj4qZMxoMbFT2qdXOFNiRTrdk3W71jXrf4EW6GFjdMFxjs02aNuknMAliFynFEuVHaZhc0jxhes6QK6hJpw0OfPo/yyx/eP0vW2pgrWhSFK7BpFnxZe1BokOykVnXKaTqnfY2VcvChG2GdVqljzg68fWqd65rdsdWrtmjqVg2H8UyEXM+Wcq7FUDGhKlp2rKvVHpTBqjTczX4ZUrPgn/dvoacQj0gTsBiSbLykTkKg2Thm+jauhHGdVqt3tCViKo7Hu2q1pifTj6cJ2V4ASAnXt2RO1tDNcDKNzRtN4ZsLnh2fhU9BwKOyI9HE+Se7Jn5+nH04W8GnLXHSrGJU+HQ6/H7Uxuuf4CEiKHyPeYom1TZOXC9LQDEaLbDSldPl2Z8Zq4zE0cx3yvi1dZpPtOh9OEYzBhOblk7OtrQj4Z6Eq9f2DdLOnmGg56Lrz0V7FFexTULFPnL+PANWwrMxPFE4hE5fOTlSZ2WrowrVwRHaLHTNC0a9A5PYEvYGnNBQPBNZF07OY2dReGXkaU6sI/WbuNpS9/VLyY/kcr1bVmCcpExiKBishXLDLSszOSrctwH7191Rpm9THM9YzJ1r9/PoPKMQt1FaPGsGkCUh0Y3RxgTVUS63Nt7nmgbUdTJrOxfuHM/bWKN3WHZeCtwZ1fYk6FR3JXTq5L7joaOfO9TCHWAPUDfdqJrchWIaClGxy0bC4sowzzjlWGtNW/wBGPM8J8fj+/wBdjQJdkOoOQTALm23hZKvBYTDsrx2V47CAS2CWoO51FZ4JXO54dVys6z9dgr6Fr1BvX2cWznH8dteK0nDZQntBkGpc0UfvTbL0iZlvRg9G7QutJqtvyfwOy2TS0bdavEQtz45Kw5KJRv4SQQRlsKQ2AD8xVgMbIc+4TEv3G+36GZsSG1c8Dw4+nCNUr6W9n4dXOdordozZ6Fwd+rx9OFZtDqQ1dOdqXeJLNcc9e6MauWvRRtcE2e8N17sF7sXWPjQeD/lbWf7tXF0fuFREIwoFK5Z8cq7a8UDXH9rKz53iyv26aLctll57S9i4vYupjXl8epGukaH4+Q13BHL0h6NbQsdnf8L8SUpSCr163Kxoz9YVevaqrveXe+u99dr6FLS507pyjw6N2Z7MvKXVqydZ9uN2twv7rQMStWxAzkjT9ha4vGAQLYovC6ojuoYNOSiPZZiexauCrbHHrbSeBh19SvJlRtRuV3/C0ISlfutLywbiNt/uV+cP5QatpRp3k1K/zcrWREFRuzZ828jZ1llKoVljBlDQvjkGTTHardJHoZPPqP8AlaNpqlbIq+MQod5TyCwlYy5uKkztM2XKKnT4f1V6q9ZTG9aVjpMcotYOKbGi64WhbapWyKzpor5BRa5WB/NaVSEX9eC9ca9ca9car1wEeyNqNnEv9HHHszuybnmnY80N3TbLpfFZNNuFaqwtB0sM1E/punqJ6rIYWjKrRrLRA1hZhYnFnWXg9O43Fa15Fwv7LX0I51TDzpVhRinZbXxwGmrecCkVx1FXhmu/u0K4G/aGnS9sVcvnr5ljlqtyYJ0dCFlvocMR2kynHs0H+warfS5fhUjcuztEvn6RFGdmdOpGuG21kMCaep1ezou/saS8+m6xM4vj/v8AQnDNcuvmaoLcDVzmc0vw6tF8K1Lv61AyuHnTu0onJpmfx6K8WivDor19J1n5+jatABEA1tWvaJQtyw7zP3XPCkLstOVqYa8pjhXqmvO4Ljv6ttercXqW16Vt01W5WjJp2z4lA2bWZkWPZhE+03+eWdozW885N19fMywu8tYXnutSkvSmo0ZoeWXgmecAatP2bEMafEcV3c8ekpx7NVn9r0Hf8XIf/KF/mXNO41Othg8YT8OKFKo6ahRTZ9Dk1SqIo6NSb/bM9Fz6DKVWqypQrhuFg3anL0rQOXWRCI5O6sP9x0hx6tz1fSzsyNn08h08QBterndJhoLxU146acdVdKqwSwKzckfLLWGuWZnVsn3LQAPqzKUfzr0Y5t2Makh/0K/ol/Qr+iX9Gm+2TrDI455tz2gs0YNzyoE9d9G8+5p1GcT0bbWRutPNFp1r2MLPN61NOCmvHUQo0ewpZIRaIWkoGaBKx1UuM8atnurJo1hVrX3zWE34+jstLIBpR1KIcsvsVEC7Rg/3uhEVecbYtmr0nVP4zVyd4jm43o6vLewNWYf1Dx4+n/1vxCan8c3ZkJf1WAxjyO5p9I2y+Unx+nxC5VtzCSWsnBpOvX0U1XSd8PHLXGmUn4a9c8qtAYo8jRnSnGbcWJtBrlnurZvMXIxykonq23f7edfbTr7adfbDIeOcksbM+3VVp2/HHqr1VrAsTRd2aTOiy8MbVUsrWqdpk+3NBvQZehFehBfb4KGWOb3hxpNlZcLxfA1QSdloVmsCxNB5Rn1nGcI3dOy0dS9ywAyr1yT9OovTqIdGi6jmZqtUaVUdCpSMmzcdU8rIJZM/YvC0qnsgyNH2AkhF9iTRe75PueiGLNA/X1xtlpo4yZsTkzZbIUctdcNT+y8TfOXakzzk01p15FHn2mtTH4x6updapVya3hCydlpNS9R7OOrxKLvXLS8RT5qc1JeaonNUXlrIVsdaxqsU6DarV1WMMwdm96wMur4RRTLhX6Ub1KuWMJls1Yy9usvbrL26y9quh3a8JaRQWDZluQCViDNHszLevuMefWYAhquZwTAWNgfVbGOLVBbq1aRu1FPOkvJUVe3RHKxo5hKs26vn2eEEjxetc5bf153FSrsAefe5TfThOytVB2obVKWZJ76DrOGT/IfKOH/yVYwpALm2+EKfZo/heR1Yb+oduVNvzav+KJnebvSHGxOTzRH4WhY4auF7Bz5pp1i07y+3WnX2uy6jjWZywsOWfD+6Zk/4V235FJlNlsAdYV+ZwW7HlfSs8RoVfdtnyhhX20a+2CX2wK+2V02VWXxr4/Cj9LdlqopScs3ZTZaQ5ALl34aINRq9yMeMyjSAM7+lUXo016NJelRTUqC9DP8AEWUSm+P5VLj+7p2RYrQhKoeemEufUkOkPDqQmPZOMdLx0V489dM9DHmKAsZXo0gxpfaWg08FZDZJLKZuUSCv9865SMOxoadj+oz63riZuI2JNCsO5nRTaOUo6WVzYv5s0O3nhX3PIU9PKRbtF39qoqpYnoEj2i7jzdO8YYLUzfdNEUeGZf8A1Hp4n2s9XNKiYWZaHAhNqlJp6Vd174F7wU9wSe2NY90ps1688o9baDOUZy09AMeGj9eF8lpsEwLsYi+4MvuDL7gy95e8paHcDO45ZN9oPauQphq9rtoUFFMqVp6xYyacXZbeILSgaVauX2qi9usvcrqrrVgrXt170oS6Sp2O8RTeL+oMphR4TMqN7hf3XH0dkQTTbdzTU2e5ZQtG2J237pIaYTzQp+OdKxyw58tyrH+d/wANas9nL+EabMv7vJWidY2CeWeRmNcFLKkvtC+zsh4XklhfH45bf3XC/srlvuuqeCJBEr+dS6AHZL0gYnlnm1KpwfbaS+20V9uoL7fnr7fmrE+NVTmaLQjMrDjbsStlZlwiRVqDPGvPwXRZtcp9O57lkIaDi8GavDmLxZiYWYoByOdNqwJUIVSEhUDQrLj6Tj2V4PMRNBjzryBOvAcVv2q0rTEoLy56YudyOxkso2cRXZg9ivfyoR+6Y6yrFE9d0ynwtiMfX+PP1IIcSaITDXki6tEYVYetWio71Rk3yGoyt7lWwOtoV6a+/wBNPvVETWrzT6IVk2oWMx7Q+NTx2YXW4ysgowxhfEy+4AZPqAVXWF7N/fHTtv8AJwvEtiJbDb7ihPbeafUdfcpJ9CTr3pKjqOG/oZcrD6dqQ6mRMcRjlFOeDL3AxX3EC+5AXtVrsJxJTsz1yOz6RnX3Ey+4GXvGXvlRyuctMvSYOujUqDas412jFeeC9obLP3gVnf5DRQTQsi3cSB2ldrQf7hXX3AC+4iUdqEQqh27BnyhyeLjm01HhdmVLQ6P5Iuu8fo7KUFt5RPG9i8yjcvQV/XtHrLNjJxBf8d0b/Nb/AMLqx/ql/r/+pq9/oVT+zp06+Lf+y/8Ar6G/x/8A39Cf2b/Q6v8A+P8Aj+M/+sktD/xmTJ/pc/sf/NU/9Qn/AIrH9g/5T/5Pq60P9EP/AC7H/h4/+bY/9mm/gMo/2Xx3/wACX0sf2u/3zf8AIf8Ayw/1U0X/AMRvrY/tH/W30f6V/wD1Q/71P/Kuf4Kqn/cKGof5NT/y5q5/kp/6XT/SSmj/AOfR/wDW2v8ABl/3L/Z/7wUUyj/r+Sf+0of4/rJWPoD/ACUP8mh/5/8A9T+k/oL+2H/4Ev8ATp/+c31tf41nf5BKH9q3+Un92TJv7C/vH/SnUlsf+fP/AET+lb+1b/Cv/8QAOhEAAgIABQMDAgUDBAIBBAMAAAECEQMQEiExIEFREyJSMmEEIzBCcUBicBQzgYJQkaEkYGPwU3Lh/9oACAEDAQE/AZSdmp+TVLyapeTVLyapeTVLyapeTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5+TXLya5eTXLya5eTXPya5+TXPyepLyepPya5eTXLya5+TXPya5+T1J+T1J+T1J+T1J+T1J+TXPyepPya5+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+T1J+TXPya5+T1J+T1J+T1J+TXLya5eT1J+T1JeTXLya5eTXPya5eTXLya5+TXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLya5eTXLyapeTVLyapeTVLyan5NT8lslz/AIhlz/iGXP8AiGXP+IZc/wCIZc/4hlz/AECH/hCXP9C/8IS5/oF/hGXP9C/8IS5/XrJ/4Qlz+ss3/hCXP9C/8IS5/oEP/CEuf8Qy5/oEspf4Plz/AEUv8Hy5/on/AIPlz/iF8/0T/wAHvn+gX+EXz/Rv/Bz5/o3/AIOfP+IXz/iF8/4hfP8ATP8AwW+f6Nf4OfP9PX+Cnz/Rrpa/8lqSPUieqPFfA5yHY5NHqSR6rFio9SJa/wDsx8/1LX/i9SR6sT1l2HjM1yLby4OBeTuMYmLk4Ocro1yQsVnreT1YmuJf/wBivn+pf/hXKK5HjRPWPXfYeJItvL+S/BwfyXfBwLyPxkiXGXDGJnGVnGV+ctjg1PyerJHrM9aJ6sWWv/Pvn/zDnFDxoD/EIePJ8DxJeS28v4P5Nzg5LoryWUc7I4OclvvlElxk/OXDy4KLKL7MquMtzk36dT7CxJoWMz1vsetAU4vv/wCZfP8ATrJj/qHOK5Y8eCP9R4Q8eQ8WT7m75ZtnubG5sjdmyLs2Rdi2LvgWxd7IWw32FsSeUuBD4FwMTtDE+2SfbK65yujk4OTctPK8ryvo3QsSS7nrSF+I8oWPFixIvuWn/wCSfP8AVP8AonOK5Y8eCH+I8IePN8DxJvuW2UbG5sbleT+CvJa7FM4N2VRfgobKvnL6sm+yFsN0R85Ld3lLOPGS2dZS23yasTOS6y44LsovzlwbM3LKLNjctZfyfxltmpPsxYsxfiH3QvxC7ixoMUk+/wD4x8/1Cyl+o5xXLHjwR/qV2Q/xE3wh4s33Lb5ZRsWz+S12NzYvxlsblJF+CvJaRuyqGyr5yu+BJIboq+cm+yEqyXud5SdISpZfuzjxlLZ3mtnWTXcTvL6cmi/OXHBeV0cleC/JybmxWW2V5b579FtdxYk13PWmL8T5QseDFiQfctP/AMK+f6p9TnFcsePBD/Ersh/iJvsPFxH3Lk+TSbI3P5NuxufyfwbmyL8G5si/BXktIt9ii6N2UN0bvnJsrzk34EvOTfZCVZP3Os/qlnHlvOHGUt0J2spKy7ye25eX05cm8cnubrKi2ucq8F+TkrwXRs8rNnlfnLcs2ZvnvlsVkpyXDFjTQvxD7oX4iPcWPB9zVF8f175/qbHOC5ZL8RBD/FLsh/iZdkeriSN3yz2n8G5sX4NzYvwbmxq8G5sajc2L8G5VFm7KSGzdlF0bvO74Eqyu9kJVk32QlWUn4Eqyk9iO2VkOM4vNeM+HnxnxwXeVVwJ3lXgUvOVF+cqN1yXZRuWUbllG5Zsyi2bFG5ay3z3y2ZRckLFmu4vxEj/U+UL8RAWLB9y0/wCofP8ASOcV3H+Igu4/xS7If4mfZDxsXyNt8soo2Rfg3KXctdi2UWkW8tkavBuykjUbsos3Zp85avBu+cnKjdlJFmq+BLJyoq+cmzeWbfZCVZN0Lzny85cCzjm+c2rE7z4zaLyaLrnPdCeWnwX5z3RZRXgvKjdF2Ubl5UbllZWc5WXnZs89j+GKU13PWxEL8S+6F+JiLGg+5qT/AKJ8/ra4ruPHgh/il2R683wh4mJ5HqfLNKNstzYs3K+5aRqN/JSNRbP+TZGrwblI1FsrycF+Cn3EkN0avBXnJyRuykstXgq+cm6LcuBJLJyoq/qzb7ISrPnNsWcuhcvNieb236F0J58ZtF1znXgvzkzc1ZUboTyouiyjcsuyjcs5KNyyjc3LKNyy0yjcstZUapIWNPyL8RIX4ld0LHgxYkX3/UfPXY8SK7j/ABGGu4/xS7If4mfZDxcR9xtvlmkSKExt+Cn3KRfg3KOCzcrycFm5RdGrwU2VQ2W2Uzgbo9zNPnJuj3M05OVHuYlWTlRTlyVk5UVfObYo93m2+wlWbFm930d+hc9C8f0F51XBedeC/OVLK8mkzgvyWjbK/JZSyvyWillZaKWextlZtnZaKWdo2Kz1MWJNdxY8xfifIvxERY0H3NSfS+Sx4kV3H+Jgh/ivCH+Jm+B4s33N3yykbG5X3KiWuxbP+TY1IbZRSLRZRSLRZ/JSLSL8ZUjYvLY2L8Gm+RJGw2imxJI2G4o3kJJGw2kbsSSytIvVwJJZbF3wJJZ34F+gsqyXR+79B/0PBfRedeC89Pg3E8qNy8qNy8qNy2WVZRuWclG5bOTSUzcsoo3LNijfpUpLuLGmj/UM/wBQYmLPW1ZbfJRSNi/sblGyNRbOeTZGpFvwblItI1fY3KODWWystRqNzgs1G7yscj3M0+crNd8FN8nBbHOj3SEqyujU5cCj5N8nIpv6s7LchbG+TYlRub5Loe/Suj9xvmzfpv8AQv8AQrOiiq46KN1znRuXlRp8G5zlRuX5yoo3LWVIostFIo3LNjbO0bFLO0Uis9jYxH72Wz3FFpGrwXIplUai2z3FHBqLkUxKhyo1HuKyci2ymyqNzUe5lZ23waW+RRo3G6Lk+DT5y3HKj3MUaz1eDTfObdFuXAlWbdFXz0WV+qxdD5yrNZ0V/WV00XQqeVIovybZUmU0X5NjYpZWu5sbFLK0bFIrK0WjbO0bFLKyzbLEfvZqZ7jSyqNRqY9RTy1Gps9zKy1Gpm5Ruai5FPLcci5M0+c9R7mKOW450e5ijRubjlR7pCVZbjlRTl9RVG+TZpb5KzbK/Tr9KsqO/wCvz089PP6e2ddNG5azpG6LzaTODV5LRsUsrNsqWVlo2KWdrKkVlZsUjYxPrZZqNymUWaj3FMotmo9xpfcSNzUe5jT7lUblltlN8lUbllt8GhvkSo3NzX4NMnyKNcG5uOdFSlyJVwbm45Ue6Qo0bm+W7Eqy3y3K6a/oa6q6a/Qe/TznRWVFFFZUiiiiiiiiiis6KNJ/JsUUaTdFooo0plMvybFGk05WsqKNy86WVlrKkUUzE+tmyLNSNTN2bFmo1+C5GxZqNZbZ/ItjUORq8G75KRZZqPcxRLLHKuTU39Jpvk4LLHM9z5FsWWOVFuXAlRbLLNRXksvKzd57m/Rv+jvlub9bz36N/wBGx+V03ezKrpq+P166qKedFFG6E1lRpRTL8mzKKNJui89KKNzbKkaSmcFoxJe9m5pzbRfgq+Slm5G7NPk2ys1eDdlLNySNTfAo+TZFosc0i3L7CUUWiy0Ofg3fIqRaLRY5eCl3ystFlmxZaLReVlllouyyyyyz7lllllnBZZZZZZZZZY9yyyyy8rLLzfnpToarjpvsxquiy75OP6eyy8qytl51lfRpNyxZ6T3F+c9ya97KLRTZp8mlFFI2KZoNKKKLXYps0lFDRqXY0tigllRsOS7FSfIopcFFZOS7FN8iSXRaNN89N/0XP9E/1EcbdKfkarpT8jVdK+5Xjqrx/R2WbdFlmxsNLLV5LLLKRujV5LLRY6Z/BcjEvWzSbm5uaj3Mo3LZbNR7maH3KaNzcbaPczQ39RTRublmpvgcHLk0tG5ubjm+EaXLkqjc3Nxsps0tG5ubm4t89+iiiiiisq6KH4RWVZ8LpoXcoorporOiXOVFZUP3LqT/AGsqulOhx8dKdFJlFdHPJWVdVFFIor9DYrKjSU10UUbl+TbKhxTNHg3Rqzn9TLo1+D3M0rockjd8Ch5Eks7NfgqT5FFLockjVKXB6a79Ln4Kb5FSzss3Ykl0t/rX02fSupbsu8rLLLO3XxnefK6uCUWjcplMplMS1bGmXgplM0y8FMVo0/E0S8GlmlmllMX3NL4Keelm5pvg0M0soo0PkplGmT4Ka5zaa5Kso0M0mk0jg0UyinlRosaKNJpz0WLYWV0aikzT3RuYkXqZos9Nmhj2KNDHFijKzSymhsSNLHHyRspm5eVMaoVlZJ+ctJVHYrJbc5UUdqKKFssqNI64RRQtMUd7yUbJU+MuT2xSLyh5ZJ6neSVjaW9Ft5YdL3MbyjySktOy5zg4xW+cHTtkp3GiyxYlR05wnp5JT1JFlnqXHQWWQxGtic3Lct5Snrj/AAb5Qm2tJN29RZbRJ+otWccS9iS75JtboklP3LNYjezHGsk3HgdS3WS2NV7McayTaOeM+ec02j+M3vycF3lwWsqLNVjimbo1IocC2uTUmaUU0X5NI4+C5IU0ykymi/JSZofYuURTTNSJJamOcUapS4QsNv6maYxL8FNmlIckjU5cGi+SkjV4N3yKKHJI1N8Hp3yJJDkjdipDY2xRKobo3ZSRsXfAlnycZc/ofT0XklYvahu+corUSle2aSjsSdu8uST7ZxRJ2834z7D5z56I5981syuUVkh7Zbp2bP8A5NLWUW0yca3z1WaHexQrQ42tSyoUvJV7ocWuSmVqKZQpVyXbNLq86ebfgh73SyrPg27CkSTiVZTRybDoUiMXNWh/cp9jcvyOi2uBSvYkmuSvBbXJY6N+wpsW6KN8npZUTFXuZpaNUha2aWuR2u+T3NJckJyZobKfkqnuPc0m4pS4NDZoruaPI3GqRRRbQk2en9zTeyKjD6h7nGUdxxHFeRYd7knHiJWdGkUdTpHtwlT56Irux75YeHfuZiSXbNW3Q32WVNuilhqiUreVkfbG88GKfuZN0v5zjyc5MdWl0d80Rqnmy806qRiKpZWx/TecHvQ16ka7rOLv2sdp088LEMXDr3LgRbRNalqWak0JxxlTJRcHvldqmPbOGK47PgcFL3QzlHxnbW6FiRltMlBx37HI42NVnHEkhaZ8bG65KHDxnuuBYvaZs/oZdcnpp8DjKOabQpRfImVGQ8J9jjnKhTaFJGo0xfB6ZOLcmemlyWo8Dk30xg5GiMeRzG76N3wRw/J7YjZqrg55zjCUuBYaRKSQ/wC41vt0KDfJsuC72Q6hzySm5c58iVFiTkPEUPbDoS85WQh+6RiYjfRxnBLDWpk5ZpWN3luyWyUCe7z7ZpWzlvoXPRH7FZPjoS2aPrimU8l46FPTTJw3tFZP3LNX2I4qWzJYbT2KFsSjfuWatCxIy9syUHF0UfyNVmtSdo1xnzyU8nGyqzi5R4HOLFbH4Y4eDjNSkuTWuxGWokl3NPjo1NcnqeCM9WxKPkrx0a65PV8HqKezJQ75WXlqo1olNqTSJW+WWzWcjN3waa+rY11tE3ZbLFcuB2hCjLvsNqO0Wc7ls1C34GnwcCU5csk4x2iyi2WLfZDTuiMWhRciahFUXZZYlq4NNCixQ1DhhwW45XmlfBo08lMSs0RhHcnPWW8ktTo06c4QSjcjEnqZZYknsSjo9ueEqjbMRlvKkySp1nh8NnbPYrd9EVTz2KVZWJ0yC0y0j9rrLbuSitOssvLBl2MSLi7LFSJQWnWiy28sHF7MxMN/UhMTSHCNakajnLCxq2kThr3Rw6YjQmriW8qIYjgJxxkSTjzloTWw281Jw3RHFWJtMeE47rKotD1LbNbboWNe0zQpbwP5Pa1Q1Jc9CxZIWif2JQlEtVVDvojOUeDXCX1I9PvF2Wkqa6MR+99Eb7HtXJrfbbqUu0TRW8j1FHaCG3LnoUfIpdoiTfB7MPndkpykV0YcW+DaPBS5mSxb2XQlZHbg2iRg588EsSOHtEbb5z5F7OMt5OkKMcJE5ub6Ir09++eDh/uZjYn7V0Yft94227eUY65UTde1EnbzhzZd75r24ZLhLoTvoX1dC7ro1cSMZb3nF/sZxnCVFLEiVWzyhLSzEjpfRg4urZmLh17llFuPBOF+6PRhYzhsySjiq0NOOzF5RJKX8nHOabjuiGOpbSHCt4lolv8AUOLXRDFlA1Rxf5GvI1SNPjo3XAsW9plJ/Sy2ilIarOiM5RNcZcjjWVPo44NT7nteeJ9bKosTRu+hJsUSSaLNdKon89FCj4JQa5E1Ec9RVdMYOXBJtfY9WuB+7c4zryMUJNbFKG8z1m9ir4zSsW3GXpyasbjgoeJq+orxnFafcx75LB7sxMTQqRalyVlFanRJ+Cj7EILDJz7mzKeXEcv5IJSekxdtkSkbPg4yic5Lc/cSpOivGX7sqNkJ6lRGsSNMlzTKvgZLdastPktLgwcTehwUnZ9mafAvctDGtLpiVlJcmprgwsXVsz01W2STW6JQv3LKi4o9SRDEWKqkemq2OHTKvZji45V5LS4FOSdkZxxOSWHa2OBwvgewk2bLk1PsKTiQlBvclhJ/SSjW0hweVFpFsTow5w4Z6af0koIlFxy/kcl2Hb5E6I4mHw0emp7xZLDaOOcnsN+M8TFqTUUNylyUNG64NXk07WRjZpUfqZLGraA25clDys9Ot2LxEWGlvMlj6doFuXOdsXudEoaeTngjhVvInjVtEbcnuVlZCPqcFKJu3sQwq3kYmLpG3LfO2Qw9asbS2R/JDDb3ZiT0Ib1O3nq8kcNVrY5W7GzDhfuZOWlDep3nqvkr01/OeDG3qJPsSdvK6F7nTRKtVeC8sJb2fVIfOVtHJHjNFbk+crJ9mh7M5yi/cQWmWkxo1vlZBJvSN9s06ZhvUjFg/qWVmn1Y33LbzTrcw5+oieHq3RfkjNxJwuOvDOec+ODCxtW0iWGpkoyw3uKfZmJDbVDpw8ZrZjhHFRPDlhkZqT9xiYb5jx0xxHEjKOJsSwXHeBGS/eTw2t+emM5R4IY0Z7TJYdK4MuLVPYlhNdKbW6Ifie0yWjmLHU1vsODXRNe9ll5UR+x95Dx3VRN3uysryUG9zUo/SKMpfWPGjBVElKU+SuhQvk16dokYOe7NUMFE8WUyuiML3Y8SvbEjFzIRjhoxMe9o9MIXvLgliXtHjLCwq90jFxFBDbk7fRhwv3S4Jz15YcPUe/BL2mJPW+jCjvqZKTk7eXLorQqJy2vohs7FvvkzC2hYnz0eRZo7ku2chu9+hviRJa45/cxN/d0YUmmKmYkNDyTcXaMWN++PRGTi7RhzUlZi4evdHcU3AnBS98OnBx62kNxmqJ4egUmt0OKnvHphiSg9iOPGa3JYXeJFywxxWJvEaa56OCH4iS2ZN4c+RxlDdDqQ010URnKPBrjPaRw9mOnyaepSou+C1wyr4yxX72WRw5PcexYpXwVZWV5Lfg9NpXRu+T1FHhDk5ldCTfAkl9yUJvkqOHyPGY1e+V5c8Cjp5KlPgWA73JTjhqkPE17M010Rh+6RKWojhSktiGHp3ZiYunZF6yqzhHWTlftQth4La3FtsYuLvRSfGdXsS29iy70hYeh2Ykuw53sab4z4jWVeSNSeknUY6UKq3NV8jWT4Flt3E7ux/Ufss2lyNUMXGSVm0eBPVEw3sYiUd4mz4yW9xz0pfUavBhTvYaUuTEWjdcG0uCMtLpk46HklfBaia5XZh4mtGiL3Zix088EXp3iTgpLXHNR7s1V9JCbi7IzU0aItUSjpe41r5GtLp50o/UOVkMRwE44g8KL+nYlFpe8lh1us1uakvpyjiOJCUG7PTjL6SeFKHPRXkcq+nJTaMLEglRLBjibwJQlD6ujj6hyfbLUep9h4TnNn5eCSxpS2yo0mtrku+M4YDe8huOGqiTxWzdlFGrzlyaPJHDvnYtQ4J418HOXBafI0Rg5D0w2RDC7zLoxMbtE5yto2kUyMKWqRKVsw8O/dIbMTFrZZUamjaXBGLk6JbLSWYUP3MsxcSlSz1dmab+khFwWrucbs5MJfuLMR7XnqT+o0N8FapGyGzBW9mJuSVZLY2fJNNIryX4yQ0L6XknRSfAovdGyG7yw3TI+xklqWSY/MScf3djV4zhKmJjWpUNU6NV8iqcdJKOjaQ5N5wlodkZKSsaT2ZOLgyGITwlPeJajwc85xk47ow8RTOVTJReHwKUZqmPCpXZq7R6E2uCGNfIpDw/3YZKKl9mSho5HcumOM1yQxVLZk/wAOnvE0b0yXsdHO76Y4kokMeOJtIxPwy5iVXJq8Z0VljYz1NLKuhn8CV8kYww1ZiY98FtlFZNjMPDfL4NWqVQI4aiYmIkSk5dWFh6fdIbcnpiQwVHfuSajyYmK5bLppvgjH0o+57kpOTMLA/dIdGLiVsuhkYObpE2sOOlDdmFh63bNkTmoobt9GFDXIxZXLbKtWyEklRKuDEdvowtrkLJmGqibOXBic9D46FlHh9Ea1V0Ik7piZNVLJifqQcfHThTFIxoalayXJiJY0NS56cPE0MjKyUNapk4PDdGHPRuYuGprXDpTcd0YWNq2ZyYuBXuiYeMl7WYmF+6HVh48ockMRSWxjR1oU6Wmasnhd4dSbjwYf4rtIxPfuh2afHTWUMecdhSjJ7jw1yhqunEXved50aTXQ25FFZWWJN8G0f5NMp7yPbAnjN8dVWLTh79z3YpFaOCeNpJzc3v0pNuhJYK+425OzDw0t2azGxuy6eeBVgx+5u9yMdTI1FUSZiSbfS/y46cku5gL9xJm9NrpltFRFk0x7IjyNN9D7dGlokIUXm9mmPnNJvgjvCiBjK42U0Mi9MrMRVLoiq9xCRqMWHu2NPdEJ6WYsf3Lpw5+n9RrTJpTVGhrYg9G6JwUlrh0r7EcbRtI1WYmEpbohrRKCnvHqhaftPXp0x6ZocXD6T03iLUl1wcuw8ZSZSlvE34aPQZ9uqLPUt7CqRT7DwpJFS8GJ9bLLI4MnuyeGo99zZcmo1dmUVlZeWHgv6pGJFOqKjDkliXsjV5NPddNWYeC19Q8KN7DelE8RyE+zHHv0Ri5cH0bR5I4De8jRFO0N0YmJqFLtIquiK9NX3H5kQw19UykuCzEnqNV7SHGs8NV72N3uKNbyMP3PcVIm74MR9kXq+oaaySt0PdiLrgwqptkxcEnxRakNVzk+VklZengT7DF/+7E37rNpD25JDyUb3Y32QpaqFsxMxtpakbTX3GfXCvGdKPI23yYchMWxix/fE2nwQde2ROOl1lzwbQ/nLCxNOzLE6J4alvHki6exOF+6OaVlpfTlDFcCMtSsTocFLeHJKOrZ8jVOs0rHLtHKM3EjiKYm48E8OGP/ACThLDdS6Eu7HK+OMk2uBTUtmRxXH+B4cMZWieHKHRst5DerNToh+I7SPVgYj97FDUyGEobsni+ByvKihe0u+CxsjBzIYUcJWyU3L+B4ijtEbb5yo3XB9XBeUIOb2IYccJD35JTUSUnLNNorVxlCDkRV+2BGCw0NjdGJiasqE9JSl9OUIafcyUjCh+5m5uYs+2ak0NXvES1OiW/sRaibyZGOlUOy6Wp5qVbMce6I7JyIxHLsh7IhtElz/wD6dqHzlfZjjW6G9xLuy8lyPKXOWrtImqRzFFaeRtvKPBLfcjRiK0MUr2kL2Oxx91I2jxnwQewssSOl7CeraQ46lTNLZqraPRhYnZ5IxIa91yQn2kYmH3RXkbvZFZwm4cEJ6zcaWJsyScfZMlhtcFafqG3LphjfI54FWIqkYn4dw3iJNm0eT6t2V0Kco8EMW3YqxFuYmBQ04lqJyV02yUbmyo4StmJjOXGdZsYrkQwrYoKC2Jz33JTb6WMjTVyMPD1sUVBbDRPErZD36oRco6pIgvU2jsKOhVEoexiT1dDyjh+zVJE59jCwnPc0lGI9COei2uBx0wvuN7VlgYf7iiSMZ/tXRbXBjbVEbsXJy0jSNUzE2fRbXA4/mHe84K2NbFMxFVZSE2hPSq6I8mn2EEaTEjplWVuqP9zCvx04ctOwiiUFJUSTg6ZGT4MWGqGpdWFPVszY0pmNgWtUTDbezMbB1LVHqTaMOcZiUSUYyVMdYcq5RiYSn74dcJuJhyw55SXu9o+d/wBDDxfTd0LGhOJ3HBDTXXPE0zdDblzlRWbZyKHkVcEHo3ZifiG9kc9N5L7CV8mH7SWIkieLq68OCXumSnLFddjC9iLJS08k8Rz6sHD/AHyMTFIR9Ri2VIbZKWnclJydvpwYW9TJ4mt2MjHU6KpUjcut2Pd9GGrkSlrlqyXJh7zJX/8ArFyS/wD3fpu5NiziM2JfTlPJdMGrFsxV9jHjtqyRhS0uvJJaXXTCViaI0Y8FJWjghiUYsNLtdWHiKQjUYsP3IhjGLBS90c1nwYWNf1Gokr3FqwncR6cTfuNNc9SdcEPxHyH7uGSiNfocEcV92Wq2LfccfBxz04n1vpu3WSi5ciSXB/J6nxHJy6bHI0yFHwLDFGh4iWxKTlz1NmDBz3oanJ7kYVk5aeTEbf8AHVhwvclKx4UyMdKrOfv2XTVuibpaEJdkaG/pMGOlWbEv+CcdKVjjpfQtovKrFHsuSMdF6ibX2I/8GnUrRp7xFmjvlsvqPTcVqZa8lpdxe/2pjjoelksl9XQl3Yn34JveyEvv/wDBL3Rolgyh7h01qjlP3x1dCje74I++VCbTqzUWehqbZRGWpaWSi4uulflb9yGJqWX/ALHg6pbEk8H+CcL3j1LbdkMVp7id8DjY8Np+0lg2iScHUupKx4j4iQxFLZjw/sOLXJh4OuN2TwmvchPpq9hy0+2JF1yJ6uC72IYcZPclgdhxcecsT63nYouZHCS/gm09in4G4xHJvk43Qvdv0WO2YOBp3ZKSXtiKHlFUTxb4GL3cldDZg4HqO5cDlW0BRyk1ElLUJ6Rx7rojHUx//Bhwv3SHK8v/AEYk6WX1/wA9EKitQrZ/ZEWmCqJa8ja8kVqZiy1SFLsxx05z8HJejjk/DvSmxy+45ff/AOBPY1OuROhq945dyPAjjdnLtjm33Y233Yn/ACRe/LMbdilq2Y9jjNK92N2J0cruRb+5v9yMqMT8uew1a1Iw3vpGqdPJKxuz7l2tQr8M38G/gxU/rSOfdEa9Rbc9H0fzknpItSVpFfYr7Cd+2SJR9J78E8N8pdHCtnLt5QlpZFqW9DjfYi5YfCHhwxUTg4OmLfNKyUtWy4zjiaeUVGW9I0yi7TMPFWJszGwK3Rus6vZEvb7YiWanW1C27kMbszEw9StHpvwYn1sstsjC9kRisNEpOfA9l7hz8dHBdljZWowcKt2Tne0RQ8jaiiU9WdCd7M4ybMHBc3bJSr2wEqylJJWSlqzT0jXdZJWzhfYhHX7nwX9y/uX9yU9K5G7FlevnkZFamSbm6Q3WyMFV7jV9zV9xz+43ohmn2Y1RHkvUx+zKG0Rv7scvuzhdyT++V6dz6laO4uBLTuxu2LdH/s/9i47i/wCTF85J2qZNNCYle7NWrNL7MS+zEvsyvsY0NrojKia/dEnutaEtQ32WcJU9zTT4NP2K+xX2JReHIW+6MSO2pZfR/PRGWlkfcror7FfYi7WmRJek6lwTw3zlxuxvVu+iL0shJS7FfZCuHFEoxxkTw3ATErJO9kV0J0RmpdkSXijDmpLTIxcKhw8G72HttErp4NblszCxdGzNSJt65I0kY3sRioIm5Sf2HNLhD36vuOVkYmFhd2Tk+IlUTnpG76WjUuJEttkYWDqH7FSyslLSiUtT6b0iUZq0RWlciTxX9j7Jl/cv7jl9yctXQxPXtI+j2xY2o+2JFanRdbWN/c1f3EPc+TGlb6NVbdh1GPtfJSgtucoq2X92Sf3Ynbq2T2dbjESE2uB6Wr7kKq2N3zknsf8As/8AYl/Il9mYq9vDztNaZGHDUrvgbvoS+zJR+xGP9rK+xptcDWl0yLoio3oQ/iumHvjTEv7TT/aV9iWHqXAm4SocovsTj6e9dUJaWJX+00/2mn+0S1qpIkvR2luhYereh3e/UtiEtXY0/YgpReyJwU0ThvsOXZldcMWtmheY0crcxIqLoaKa/QUnE9WRKPvZwYRi4kUqY5X1spyFCiC3ylRPEXC62fUKGkwvpJV3NiUlFEpan1fYw8JYcfuNapaURjGEaQ2i15NS8mLiftXSz8PC3qZP3PUMwY6FbNa8nqLyPEXyNWiFsbvo5MX9uGh5YH1Wa0PFXkjLVLkliK7tkneUuclsmxcDyRrX3NS+4n/JGX8mI7j36MGV3Bj6IeBu49yMvsxP7Mv7GPH92StLVExV+5d+mL0ys+9H/U/6ivwY+FqWpcmHT2Zs1oZKOh0+rDnp2Z/1FfxImNbjSVmHKWC/cYsNa1x/Qw8X9tEb8Fk4zbs5OOf0IzcHaML8Qp8mMnIqlvk0fz10T+p0Ou5Kfj9ByFFvkSKl4FD+0c9PKMTE1vrvyc8EY1wRjLuhbdh79ictPYbvrw4+n7mTxW3SMKDgWx39jf7E5uPVy6JPQtCJuzDWt0y/uN/ccv7kRuT5MeXboZh/UN6m5Z4O0bsc/wC8c/7yL7uRq/vOSh85N13Fxn+01L5mr+8i6/cal8mNpx+rJZR2mNZRy4ZFp7WxNLlsTXlia8sklKNC2IshvFwK6cOVrSbLbcVeGKvB/wAGJHRK0OWpWS/MW3PXCSXJFLwX9h79iWGviRcsN+5bElq3gv0MPF07Mu+w4J/tJYb7RGn+43XBt+hDEpVJGlS3USUZt/ScbMas00c9WJLTJjbfPU3Rfku37SMMkk+UVFEpxrYbb6nsfVwU5bCjtSFFPlFJdj/gcorZold79eHT35JyS4MLDrdor+0r+0r+0e27iTVO+lujDTitbR/cxrwYcHFcG/gd+ES1fFEFpjY1qWrp+mDYhKym/pIpqNbD1/Yev7CvT2Pf9hKnUhbbHfL+cmJanRp1+2AnL5IuXyRFu37jU/mjU6+scHHdjSrUspckvIxcjKVqK5NUk95jel7SNf8A+QU/7zWvkPCc23FlWrRel2iXO2V5VbpDdOkS23TFJfI1L5GpfIemSpsUJb0RbXBNLldUV+5kMS/qZcfLLj5ZcfLJKHdswYOTdPYxVo61HUxYm9dhSi/I9P3HCH3yWHqexLC0vSz6XUutvQtKIyjVSKh2TPcuxY42SwvTp8oxIV7o8Cec372n1OXghDStTFhqKuYo0bCjXctLuSxG9i9I146WyMZYstIoxwUOrIxXkteS15JSS4Y3qF71T56t5vSiGHfsiShBLSz2ntPaXH7kn4Iv9suBrS66ErZSk/aV60tMeDTHDjpo28Ht8EtPxZGMZPZGJLT7aE9Lsku66JdlRzsT+ERL0o1FFf2Dj/8AjNK+BJbL2WRuLtQMWTlLcvWvvm837FXcwJSjelDTf7DS/gRT1fSaX8ELV8EO5xepEJVsxrSyQvpQ8k9KvuLZ2NSe+lElJpNoqXxQtfhHv8ITmif5eJfZklRG5Rrx0XoX3ZRhytaRalse/wCx7/se77Ccu5i4X78Mi7W3BOOl9CWok9XHGWHiSltZ7vJb8lvye6P7j24qpGJB4Mvt0/wSde1ZRlKHBGba+ot/Iab/AHjqHDMOaxFpkYuE2iq6fo37iyU5R4Zd/uKiuGJ2YeJ+2Q4aduzJwp0zdFmL9bEtX852kbsw8PUzSo+6RJ2VLsJPwSnpJScs4vszjNuitbIQWFGyTeIRjI9x7ic3Ee+f1b9Dd7Iw8KlRtFVE38m/k38lv5GJOXF5x9y0s4yYvavayXtWlcsilhR0l/3F/wBxq/uHL+8hsrkyTt85QlWz4Je3JU3ucuz6F9zDrVuNx+RcfkPT8xU+JEnD5Hs+bHycO0Pdall3yXtWrKFdy8Pyz8vyxOFn5f3F6f3PZ98o+5aRkOBiXdjdu8lorcjo4SZ7O6Py/DFo8M9ngxIpx2RB2tLPpluSWUfky9Tti3y2kroWl/tNvibfE2+JGWnZRMWPpSvsylVUU1s8uR7e1dEZKW2kr+w/6Gm/2Hug/bAlFYsKZJPClp6H7FXcSz4ZCer9pT+I4v4jhO9kYOJqWl8mNhaXaHGuM1stTN3u+mOLe1EoTfY0yitzBxL9rMXD1q8tjE+tnBdqxvwaRK3SIQUEYkxKMuSoIniJbR6ovs8pSQo3yYOH+5mJO5V2FGHg9vg9vglKK6eBruspPwfh8G/cxuh/wf8AU/6n/UlJL9udZf7i++UE/qoW35lGBHVJ4g9T7G/xPd8R6vgU5OnExG4qqyZRF6lpYzeMbIKlqY3Zgxlyke/wfmeEfm/FCU73R+b4R+Z4WcXpZNaR3e4lf8EnqeWFq/afm+UP1fKFr1cl4nyQvU+SPf8AIl9TsRJalqIeCrdEqeyzw3LhOi8S/rR7k6Uj3/M93zLl8zf5DWmVH+5H7i90d3wJW6RLwsolIi96N061H/c/7n/Y/wCwqktMmRvDl6b/AOCce7e+X0L7sXQnXBFqS3kbfI2+Q1H5EJRw39Ri4axFZ/tunkvatTOd+qEk+WezyVDyXCD1JkZLFjZOGkaFzUiT1dVCdcn5TJOK+kwcT1EYuH3RRifWxivsJUJGHCtzEdqkRjJcjk4oniuXWzUKJh4eonsqRFS7s93k93kniSj3G76WKWnZ8E04GDhOTFUUP+T/AJP+x/2G/wC4bb3fTbjuiliLWhR8PYl+ZLTE9qVJlx+R7fke35DcPkRSW7ZN29mIeTF+b/I4JyUUybvZZRUEuT8vyP0/LH6XlkVh1fY/K8sfp9uiO/sZp9+knS9qzjp/cfleBvC8Fw8F4fxPy/iJ4fxJ1ewiLpjSjiUTqHtXQqvcej4HtcbouHwLh8D2/A9vwMVd0qIOtxuCeryS9i/kWadjI+9cG3Gk/wCh/wBT/qf9TEg8aF9yOIuJcmj99G7ds46U6dkZauInu+J7viO3+0w3Jr3Ix8G90R2lUuCXue4uuGK+D3+Cp+DC9ROmticdSGhqzj9BNp2hYsnsQWJqOTQjFfvYoiQkQ+rJwjdk5RiNt/oPcjESI7InFPkqJUSbiuOvkasS1cmCqQyl4NvBt4NvBOSb26nuQw1hYds3gtR+Gw6WpjX2P+D/AKn/AFOXTiTeiPGXHR+Hh7nIS1TbQ1RBapUb+D3eB6/ifmfEheluha/iYrenddEI6pDp4xNU88C96G8QvF+xJztXyJ4v2Ln5R7vJj3avJfcxPZNbGMt76VKbX1G0o1ZGUvJcvJb+Rv5GtWzYva2jTqVodYmEnk8ousoy0sns7iy/7i/7hPzIuPkVH4mKi9aMCepUzFw9D261Jx4E0/3G3yNUfkRaoxZJR3HTdCdcnP6EJ1yXDyQcew3SJTjftebVcfo4eK4ckMSMzUia97KySb4IqS7Fsnj9kc9fB9Qo0cChJOxau5LV2PeTxZR2OemyrNhLUKF8GHqX1MZ7vJ7vJ7vkTlJbX1UYS1PcnPU67H+7OuyykvuU/kU/mNf3mFHu2YruXOUsqKHNYeGR9uGcGClJtsqPyGofIcYfM0w+RJRpe6jTD5kklw7zojSdkacyXOcdH72Vg+Wfk+WP0/2lYPln5Pln5JiaKuIssZWky1KK6Y+nXuIvBUiShe5+Sz8k/KI+mY6SepEHRCWmVPgapjzUjkw2mtLKgvqR+X8T8v4i0fE1LwYzg/qRq0u1weopR4Kyvpi0nuaofETh8RS+xOSapotL9g1aE9G36MZ6exh4ikrSHN+B/wD9Bub/AG5uPgvroVx3R60if1M4NN8s0/c+nuSm3+g2K5CVZKEe7FFeSo+So+SbS4f6HA92bCWGz2IuBeGXhknh1t1vYc4KNLklJw9hhqEUa4+Byg+w5YfgcsLwL05cIcowVUfwX04klOVJDGYVRhuhyj8Ryj8DVD4Fx7RolON04GqPwJNPhV0WYfI88NtcRs1P4GqX/wDGScnVxo1T+Bc/gKWJ8DEc3HeIspbog24V04baeyNWMuIE9e0pI1YvxLxfiXi/EXqeDEjOcaoiS8jbxI6umJ9LsdtakKWKz80XqH5g/VJwxZKmRcsJ0xqeIryo46Y4ko7IXqn5h+aP1RxxnyONOmcZMXVGcocEHOavUVifIcMX5HpS5bL3rJqzdfoUYn1sWnuewlOK7Der9ByFGxLJV3QtPxLXgteCeIuy/Rty2QlsRb+Jv8TU/Bql8Ryn8Rzkv2knqfWtcXaQ/e25GFGcnqovE8F4ngvF8DeL4NWN8TD1S3ZiSm3pZx0pSXugRtvU8vqdH5qPzj88/wDqBeo3Uh/6g/8AqPI9Upb9DvsYedWrIKe+l0acX5Dji/MlGaXulZpxfkacT5GnE+Y4TreZGLyfBh910JanSKp+00S+ZoeneVijKX7jQ/mKL+Zp/vNP9446Z0tzl0Q502Pbbp5IfU4jhvVmmPzNMfmaY/I0x+Q4Rf7iWHFfuIO9mxvS6l11ewo+7TqPTj8zRH5miPyHhwf7j04L9xsz6Wckva9L/Q9iemRWF5HHB8lYPk1LJqymuBprZjuDp9T1KTpGprlE8Vvge/u6nsJSxZUiOEpOkSw9MhIpvZCU48HvPeXMxMRy2PrV9e+JLSiOEv8Ag06Ze0UMRFYnkqfkqfkqfkaxPJJy8kvctaF0pa9iWuG1kMBKFSI4bjsmVL5GmXyHCXyHCXzNEvkaajVmI+yJe5aujgmqjaYtkTjxhksOFUzSvkOC+Z6a+Z6a+ZGK7yNEfmaIfMxWttI/d7851W5DLnYnyooxXhTe7NOF8jTg/IlHDX0s04XyNGD5NGD8iMcBdzHkpJTiS392Ua1bjzXsjq8mBJQlbJei3YvQTPZ3KwBf6c/JPyTDnhR4PxENPuiT3Skh6WtumL0rWQel2SlCa2Pylyi8HwasHwXheDVheB+j4MF4cvakYmFcdBGV7ZrOPtWoQvT/AHH5JeEasLwfkvsSlh9kJruTgsSOqI4+rD7oTrZi6Y+1ahIjJR5R6kPia4/Ac4r9hbyWzsnFY0bGvUh90boT6MSTi3ZKTkUL2sroborVyYcdMR1hqlklq4FB9maX5NP3K+5KWSel2NV0yd7GDh1ExJaVpQoKXcWGl3Kj5NMfJpj5HGHkkkuGURel78MrS6Oc+DTCW9mBDVLW+ETlGXc0w8lYfkrD8jjheTTg+TDhFO0TeFLKD0vcap1ndcktDl7CKr3GD9bnIk8OTtn5Q/RPyD8g/KSqR+QXgeB1ftIOnT7lVtlOqpkRkfatR3NeD8TXg/Ec8H4jnhte2Ip4dbxPUwviepg/E9TC7RJzjKNRRhvsVWxLaQ998ktTom7lscM9SHxPVh8CUk/dR6sPgLGj8D1Y/A9VfA9RfEjP1fa0Q2k8JkHouLXRWp0ibt0uFlhT07Eva7o9T+09R/A9R/E9R/E9SXxPUkt1EX5sb7mNHRLUhb5pn1PSOSlKkVl6kfiepH4nqL4nqf2jn/aSk5ftMLEcHTMRVU4oxcPezjoUdTJPVIWUZuHAsTElwasbwN43g0Yngsw56WSWl60YkNLKE/OeJ9bzaFuqzbKMOGtm0dyTvdi9woQ8mmJUT2+SUr4zZDdaehvsjCw9THUFZqi37hLDPYew9heGScOxWUtyHvjXddCkv3DSk9MO5ccJaS8PwaoeDVh+DVh+CU8LwXhS2US44cd0SlBr2rOPujXdZ6ox+pWQ3ZN0tKMOSjGmjXH4muPxHiQ+B6sPgepCW2keJGKpxPVj8D1Y/A53y+qP8ZTdKiIlqdE3bO48WXxPVl8R40viPFlJVpI4skqUT1ZfE9WfxFi4nxJTm1TiLgfujZMtyV5fTG/OccTErZHqY3gcsWcd0LExOEj1Mbwa8bwasbwasbwasbwfiE1WIS7YiHqmtTz+iN92JZcEZSxImrETpF45eOfnl45+eJ46luYkFiRo3i6fQ/ZH7sihPJPS7R6s3wjXieDXi+DVjeBvG8Eliz3aMCf7JE8PVEcTjJuiXtjpF0W48EHOXDNGL5Hh4vk9HEPszClftZiwuO2TjZwWYi9z6Lp2NfuRfgUcsKGlWYshNN7nsPYXEuBOV8ZvOW/uyk/AlRhQ0xMWa1UJw8GqPg1R8GqPg1rwepH4nLvJlEXpdkl3WXY9RVwfh4UvUZ6l9j1Psep9j1Pser/aPG/tIPW7onjSuqJPU7zunaJeVlKclHRRBaI2MU5LsepPwepPwPFxPB6uJ8T1Jy2aHiYq2o9XF8DxcXus4vS7GtLJ3/wR4H7VXnJXexeOX+IL/EEvXr3EXjafaX+IL/EF/iD88RF0YirYjbiJanRJ6nnhuf0wGvxAo/iO4vUT0xK/EGn8Qacc04xpxjROUWpGF3jIgp3oGqFHU6JPVK+jDk47E4tbijiSV2eni+TRi+T08XyaMXyPDxfJgqUVUz8ThfuQnWzyjG3vwiT1O81uUJuPApYsuD84rGKxhwxj0sXVqIu0Y0Kdoas+khv73wjdu2Lp4Ie/uel/cPAfyPR/uFL05EXqVmJHS8mjSif1MoeabqhLLDhbJPTETt3IuPguPg1Lwa14Jz1dcXWzJ+zYijChqZKWlWLEvsa/sa/sa/seo/B6j8EpueTddEH+1leRTcN6N8aekm9CqJrl4NcvBrn4PUxPA8XE8Hq4ndC1RjsSxMSvd0x39jKfCG5Ys9Mifggm5WjVimrFNWMa8c1/iPAniye/Jf4gv8QTeNXv6Ie5aGYlrYwl3fA93eST1KjRjmjHNH4glh49bkI4sl7T08c9PHPTxxYeN5KcZU8mtcP4MPe0j6Ifd9Cu9j0sXyeji+SUJRfJ6OJ5PRxPJ6OJ5PRxPkejifI9KfkxoaJpsk9S1LsSi1HUP2Rru+rC9/ceG7qz0X8j0X8j0X8j0n8j0n8iOE09Woa1KjEhpdCl2J+1aCs0znK3HgUcV7mjFPTxfJ6eJ5Hg4nkwYyhtIktSoktLGrHa27ZrqjT5PSh8j0YfIeFD5GC1H2WTjqQ9s5/U82VYlkkQVIxJUal4NX2NX2Nf2Jz1dHPRIS7sSshHSicmnsa5eDXI1SNczXPwPEk9sryWbFeJh6iWNL6WYGHoj9yUp3sasQ1YhqxTVijljGHql9ZiPFX0kpSl9XTLYlq0LEjyYdU75YzCjOrR+afnDWOV+IK/EGH6jX3HD8Qen+IJqcdp9HDVH4rlDdYais0raSPQxfI8DF8n+nxfJ/p8VcsWHOX0s9DF8noYvk9DE8noYnknFwluWRdOyG+NsYu8ulYMpK7P9PPyLBcY22LB172f6d/I/wBP/ceh/ceh/cej/cTwPy2YeJSowEpS3MRPVv1J0aFKOwsK+56H9x6C+R6C+R6C+R6C+RCOmNH4iFrUfS9RzvlWcZUeojk3XAsPEfc9LE8no4nk9Gfk9Cdp3l+IpZND9uaZZayooVdzRhvuelh+TDwYqVp5Y1XnL6mPKQskR5yl0YnQ+mWUOf0JfUxjyWcjB+hE/wDd/Qhy8nz0z4H/ALJAZg/QurD7543K6EfiOIkfoRLKH1dMeBdEvqzw/wDdRic9K4JGFwzv1R+kw/qML/dMbnrwvpJ89KEYv0D4IcdSEMhwPOHOX4rsLKXBHjN5LNkclljciy//xAA0EQACAgAFAwIEBgICAwEBAAAAAQIRAxASITEgQVETIjJCUmEjMEBwcYEEYlCCFDNgkXL/2gAIAQIBAT8BUVRpRpXg0rwaY+DTHwaY+DTHwaI+DRHwaY+DRHwaI+DRHwaI+DTHwaV4NMfBpj4NMfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEPBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfB6cfB6cPB6cPB6cfBoh4NEPBoh4NEPBoj4PTj4NEPBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoh4NEPBoj4NEPBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBoj4NEfBpj4NEfBoj4NMfBpj4NMfBpXg0rwaUUiPH7Qx4/aGPH7Qx4/aGPH7Qx4/aGPH7Qx4/Qr9kI8ftDHj9oY8foV+yEePzn+ya4/Qr9kI8foGL9kFx+0K4/QWWR/Y9cfol+x64/RL9j1x+0K4/RL9j1x+0K4/Rr9jlx+jX7HLj9oVx+0K4/aFcftCuP0b/Y5cfp7/AGKXH6hP/kqZoZ6YsNGlCSNKZoTPTHhmiRT/APjFx+pT/wCL0sWHI9LyLCRoRSRwc5M7CyrLnOrNMWPDR6Xg9Nml/wDwti4/Ur/hVFnpSPSZ6S7iw0Ul0c5Ucj8CzXTz0/xnyaV3PTiekekzRIpr/n1x/wAxpbFhSFgnoo0RKS6uCsqyrLjJ+MmLnJZc5ciK/MryaIjwkekelIcX/wAyuP07zX6jQ2LBkz0fIsKIsOKNkb5b5b5b58HJVZVQyu5yJdx7iyXOS5HyIeTWVd8q8ZcnBycGzOMq6KyrxlyOC8HpRPQ+48GQ4SRX/JLj9Uv0ShJnozPQ8sWDEWHBdiki8ts/4yvPnOiyi8uMq7se4lY8u2SyQ+cu2S32yQ1lzlyUWV4z4yo/nr/npcV3R6cWegux6DHhSNLX/GLj9UvzFCT7HozF/j+WejEWHBdikizfp36qLN2cFlF+MuORsqzjJLux75PbJKx5ds3zkvGf3yQ1WXJWVeMuSs+Cys6Ly3/Lo0Q8HoxY8DwejIcJLsV/wq4/VIXSotiwZsWB5YsCIsOC7FRRZubZb5/zluUbG7P5LKbysqzZFlHGSRfjKi8q7su8ltvnws3nLnJbDyWfJWXJWXJWVXlZtnWVlG6yo3RsUb5V07Zbl5OK7oeFAeAuzHgPsPCmjS1+vXH6mhQk+ERwJsX+O+4v8ddz08NGy4Rv0VluUbG5XnOjY3KLRZRsiyjgvLg5KOBvKq5G7yruxu8khu8kh75y5zlm8+Vnz1fyNZfyVledm2VmxRZsVnRusqOMtsr6t0WUmenB9h4ET/x/DHgSQ8OS7FP9QuP0miTFgzYv8Z92f+PHuelhrsUlwiyzcrybZUbFlMpZblGxZRsWUbF5V5OOMqNkWUVXJeSRfjKjjNLuxu8qH4z4Wceeh5rjNPo56rP46rKz2yssrxlZyUXlWVmxWWxRvnReVG/R/Jpg+x6UB4C7MeBIeFNdjS/0S4/O0SfYWDNn/jvuejFcsUILsKlwizfPcrybFlNlZ0bZ0cG5RSLOSiy2yivJfjKjZG+VeS/GVFVyN5JNnHGaXke+fGaHmuh5roX59dFdFZXlWdZXlWexRwWbFZ7FZbFG+WxRRZZpix4UPB6ER/477DwZocJL8xcddChJ9hYE2L/Gfdi/x492LDw0Ul2LGyynlsblGxeVGxZyUbFlFFosopItZUbI1ZVZsi8kjZDeSRaWaRfjNIbzov8AL7dD46H+krorxn/JXRWW+VG5vlRub5Ubm+VFM3yop5bFFPop5XnS7jw4MeBA/wDH+4/8eQ8KS7FNdKKFhyfYWBNi/wAZ92L/AB4LkWHBdjZcItm+Vm5TyZuUxLK2Uyiy2UyvJZbKZWW+VZb5UXXBbyplpFvJJmyN8lZwPfOqLefHI7fVXU8t8n0dv11Z/wAlZ2bZ2bFZWbFZWWikUWWbFZWbFZWWjYrKzYrKzbLcssai+x6UGegnwz0PuYeFDSmbIstm5RsWblFLLc0spG2VMr7mxeWkpZclFG2VGk2z0myLyo0+S/GajZsi7yopLkvNIuuOjjorLbq2z2Nsnltl2Njbp2Nv0tll9F9FmxWdm2d5V4yss2Kyt57m5eVG5bLKKZuW8qNzfOjctkF7UUjYs5NJsbZUUjYvKikWhsSNJsXlRSNs9JsXnSRaRd5VZSL8Z0bIbvOvJfjopIu+jj/4G8t8ty8t8reVG5uW8qNzcvKmbm5eVM3N8qKZuW8qKZuWzDXtRpNi1lRRsXlpKRsXlpNKNstjSUi0cmxRsXnRsjVmontRZtkkbIvNItLgvOi1+vsv8zjp46eCyy/yr/IrO3lWdvKjfK3lRTyt5UU8reVFM3LeVFM3N8ofCijSbF5UUbF56TYvwXlRsWuxd5UUi0WbFFJcmpdi7z0+S0uC7y2NJsi7NjYSs2Q3ZsbZbIs2Nui/01l9Fl9FlnIsrz46eC87P4LyvOyyyy87LLLyvO87LLy3LLLLy3LLLyp5WajYo3ytl5Uzctl5Q+BG5RpZpWW5RRp8m2VFGllLOhRNJt2yoo0mxeemzSlyX4zo0my4OSiiiki8qKK6a/I2NjbLnLbLYZsbGxsbC/J2yXS+jYdMXh9PG6LXTdc/pb6bLy3LLLLR/GVlmo2KeeplmxvlZqLzw17EbFm+VMrzlbzpmyL6NJsW8qKZVclvsbvKmaWyki2UUUKJxwblFFFeTfsUUUVluUUUVlRRRWVFFFFHOxRRRRQt9yiiislwUUUUcFFFFFHcoroXjpasTvYrKsmu6FvlWdVwc50V1V+dWdmxRWdmxXRZsVnZZsV0QftRbNzY1eDUWWUzY1FlllMtGosvKmWkOTeV5JPuWkNt89FF1wX0UX4/RLpewlXS+p/mPqYt+lq+BO+lruJ300X56r8/o6K6KKKKNzfLSUUUW8tJRRRvlsYenSjUststJ7UXlsbGk9qNSLRsbCVj0o1LtlsbFGlLk1JcFo2NjYUV3LS4LRsbG2WyLNjY2NvybLLLLF02R8vovLl2WX0MssvN8Z3leUX2yssssXteV9DXdF2WWWWNWKXZ9LVm8Syyy8v4FIv8iy/ya6LNRaZXRZsV4HeVilRq8mxWcPhRRp8myL6KZsjV4LvOjT5LS4HJ9CTZSXJq8dOnyXXBz0UcF9KX5t11/E+qToSpdXzdTFv1WlLqe6IzT5zs1Isb07mqPktFotItDpilWzNcfJaLRaRsccGpVZqWepHJdGpGpFlmtXWVjklyJp8Z2uMrNaRqTLLNSZtlazuhSsvLUs9VGxtnWWrKElpRqNZrWVmtGockakallZqExmovKzUWNmosbfYTNRqLdmosbb4NyzUb8mo1GpvgTLHMjfLLNVFyk9srJTrZEbXJY3QtUmVlNv4YkVpWUnSIqUtrEqyxLl7UJVlN7EIu93xnPVJ0s8RXGkQhvebw7lqzxIaiENN5+nUtWeJBPcw46fbmo6JfzniQp6jD+nOK9N12zxMOtyEr2ya1bMX4ez4zlh1uiM7yaUuRXHZ5cjhW6FPJqzdZ1XAnk1Zus6rjNrorxnZsUWWUUWbMosspMplstFeC2jV5KTNLKZFvShRbKS5NdcFtlFotiTKS5NXgtso2LZRRqLK/J3y4626KvnO74EsmxJy5OMm+yFGsm6N5MSrbKUtJGNb5N0NuW5FaVWTdKyC7vOTtkFSzj5zb3I8ZrjN9HbN7oT4ebVoi7WT32N4iknlKOpUQlezzcHHgWIu+TVieh6XnKHgvTtIUk+Mn7RNPjKULEmjUrrKvApectNiiyT08iaZR/JyUaWOIpJ7dFM0mkk1HkTT4zopleRxrcjJPKhISZRoQ2o8iZsUJM3MN1FGpM0xHpRqQq8Z2bMdI1I1ItvgWxeVI1JGr7HqeBKV3IvLYdGr7Gui5YnBxnIX3NRLF7IjF8yyvOyU9KticsV2uBKs5O9kRWksxMX5YmHBvd5yaSIxrd5N6VbLeI7IR0rNrVLPHk17UYa3znwLbPdpsXVI3vrkuYmE7jmtpVniRtCfpyvtnOPzITtXni4ZhYl+2WTSZF6HpecoqQ4ywXaITU8qrdClec8JS3XIpuL0zye4nXObSezJYUo7wIzvZ5J0XecsNSPdD7iafBYpZ7PkeF9Jco/Ec8GtoUk83FM0NcH8ltHqeehwTNDOBTa5NaItKKNb7G75NPS5JGpvJIpZ8Dn4N2fwaL+ISS4zckhybEi2/hFh95dDkbj9vJ7p/wRgo8dFlEp6SOG5vVM4zbvjOc/liYeHXPRzvnN+o9KMONZydEVSyb0kd3rIKlny85OkJVXR2zY9s10T2dieiecvIt85YdmHifLLP4HmyeE+UQxbW5yNWRlWzzdPkeHKPuiRxFJbnI0KXnOSUlTFhzhxwKSOS6LzlFTFCSLXcTvgvolBMWHLuNaRPwWXm8O+BYbrccKIy8Mvo9Pwena3NDiKfYvoeGemyMU4psVIpGke3Itx7Gq/hNN/EbCSNI/byJ2Mc18pFN/EbFIob08idnI5RjwR1S5RsbFDenkTsbQ5qJDXJ2JJGxQ3p5FLUbEsRRIyxJvYjBRzbrdl6/wCDYcqNcpy2IYahm3W4nr37GxZOblLYwoaVm3Ssi9b1Z40rlSMJZvYg7V54u7SI85su10N7dFvVWclaJ7xsi7V5wbUtHRjQrcwp6lWT3RGTUtDKzx8L5kYWJWzyatUKTi9LKzxcG94kJuGzE74HuanF78dE8NTGpYLITUuMtTjzwKnnKKlySwnh7xI43ZlnuT+wmnm0nySwO8TW4fEKSZ7luRkmXm8GL4Gp4YsRSN72E+iWHGR6co/Cz1O0je7TEy8oL2rolp7nufAsNdz+Oi32HFcyHPtEWHJ/GxJR46NXgce8iUlE9+J9kRgo9Fk6XJbZcpbQIYWneXQ5UNX8RyTxNPBDCc95CSjss26Pj5ylJQQ3LEZCCh0P8V12zxsT5UYOH8z6MT3PQhKtlliS0RIK3ZFUs58UVW2b92IQ7voqlmytuhrdPolHlGBLtnNfOhO1nOOpG+HITtXlOOtGHPUt+jGwtO6MLE7SyaUuSMtPtl0YuCp8CcsJkZKeSuHAnebSlsyeA47xI4naWVd4ilfRPCjM0ywiMhUzVXPQ0nySwa3gamtpG0i3EjNPolhxkaJR4FKyzUl0Pfk0Lse5C3yjL2oTsocWUllWTkkOfgjTKPT33OOOhz8DfkU4tbGmUhYaj0Xk5qIt+D0b5EtPRd8CVDxIot4m0RYCRdZylpOd3k8VJ0Ri8Viw1D4eiT1+1CVcZSxuyMLD1u2VWcpaVZBVzk3SsnN4hhwN1nzLPEbjGzD3tsiqXQ85HYhvHN/DnuSVOyV4crRB2rzw9npysryY+HtaIzcRO8pe160RepWWbs0p8mNhad0RxWuRbjSezIy0+2WVlNmhE8N4buIsZ9xb7oqt0RneVlDhFkoSw+COLT3PiLcRO868koKROE48CxWviE73Qp+crKZSHFMxIT7GqviI4jIzUs6NkUmTw59jXKDqRHFFJPOs8PBtJyYlGPBeekc1wSmW5fCRwL+ISUeC+j1L4HtvIc72gRwG95CSjwXlyS9qsU3Lg+Hkli3tEhgXvISUeM6ROejkWqZtEni3sjDwtQko8Z0TxNDojFvdj2J4nZGHhubElFUs68EptvQiMdKyxcT5UQjrZFKKrOvAm8SV+M8afykERVLN7KyHw35zx3tRxEXGb2HnIvYwuM+zI7rOfwkt42YEr2zxPatQt1ebVmJHSzCnXteVF+lKuwlm1Zi4ehmHiadmLySgpIhPTLTM/jPkxcGt4kZuDITU1sShe6MPE30z6cTBUt0KUsJkMSMycGt4mHiriXJfRPCUyUJYTsjjKW0hxkvgIYiez26ZQjLkngSjvEU3xI90XaI4qfS0nyT/AMbvASmnUkJuDFip9EH7UUVlqJWxLshYC5kKo8F5VlLESHqlyalH4SODKe8iMIw4L6JYlcGhy3mPEUNkaZ4rIYUYF9EsTtEWH80iU1BEpSxGYWB3kcdE8SvbEhh17nzli4rlsjCw3MSUVS6MSde2PJDD0ZYuJpVIj7mYeHoXRiy+VEYqKrKT0qy9Tswo9GJutJxtkjF3lRXC6XmzsQ75oW3RXMSL0Sz52MPb29GLG0O0YU9SylHWqZhTr2S6JRUlTMTDcWYWJp2ZdkoKZhzcHpn042BfuiLVBkMRSJRUuRSeHtLgTvjonhxmtyWDKD2I4r4kOMcRGqWFs+CMlLjpn/jxe6IqceDVGfItURST6ZQjLkeHKO6OVuLUuBTXfp5HBDjQk1wKfktGH8KOB4qOTQaK5yvocqHPU6EvB6V8igol5Vk5JDk5fYjOC4LlicCwEhbbF52kOTlwXGA8ZVsQw5Yjtiw9HBd9E537YkY6SWKosniatkYeDq3YloLvPEnpIRrdjHjLhD3MLBpWy65zbpWQVvW8m6Vsnia9jDRGFIvzmt5XniPSrIe6Vs77FeM+4+c5J7UdjfXRxkuTvlZVk1plZircwZN7POWz153fBp8mNCnYm48GFLVzycGJG90Yc9ayujdjhFqjEw9DNclwYU9X8ko6uSE3B6ZZ34NN/ETw1JUSg8NnqSIyU0bw4IyUltnd8CiYmEpjjLCFiy+YjJN+whi3s87NLfJwSwlInGcTXJckMWxO87NP1ZOCZiYcrFiyw9pEMWMujng093lpNB6yjFISnikcFLfKyzTfBWTdE8fshRlickcFI2ReWnxldDxPBKfjcpy5IYHk4LOSqLJTUTee7J4naJVmHg95HBZVm6LRPEcvbEjHSjExPljlhYV7vOrN1ySmoogrepleTGn8qywcO93np8GquTElrelH8HBiy+XLCWdeBzrkjtHPHfYw9tzD3z4Iu30SLH8S6G+GcnGWIriS9yIvTLPtTMOXylec5xtDVEXpdkZWjT4JXCWojPWthKs5xU0Ti4umJ07MOamieHaI4rhtIVyFtnKKkqZiYTgLZ2iE1PZkoSg7RHFvY0+ehpS5MTArdDiKfaZGco/dEZ6+BJLo5J4KfBLCcSOM1yLE2sg9as2XHTLCUieDKG8SGO1sxTK89WFgKk2cF9LkiyTlN0YeDXJwX04mKuEVUbkSm5GHhORGCiWXnwYuLq2iKo+6RPFciKcuDDwtO76W63ZKTxZe0jFRMXG7RywsK930ymoK2QTxJamJVwYuJpVZQg5MSrboxp6YmDClvlJ6dxtt2RMONLoxt6ijjPFdyFaiYapdHfollL4l0TTq+h7iVWhowpXHJMf4c9XTjYfcaMGel08pK0YbeDLS+OnEw9aJR08ik4O0Yc1NGJh6zCxHh+yfS1Zi4GndZYWN2kTwr90TDxvln1YmAp8E8Nw5MKWlmnfVAhi9pdTSlyYn+N3iR9mzFyLE89csCEtyUHHgU2hT6YP2LpscixQEkiy+hyUeR6p/wXGHB7p7Ihgpc5X0OSQ3LE/genDJNzZDBciMFBbdLkojbxn9ilFUYmI5bI02YOD3fS3W7N8aX2NlsTnoRK5OyMbMOKiumP4ktWTfYxpX7RIjzT6Y+6TY8mxbsfAmlt0LockxExSz5iR4zuie07JowpVIsRKOqNGFLVHolvsYkaZRhYm25qMSGtGFP5X04sPU4HCiMnB2hYie5NKZh4jg9MuqWBrdxHFrkw8Rx2ZPRIjNw2YnfHTJJrc/8e90e6DE1PkWJ6b0tid9U1FrcWC0jjkXOx66E76pRFhbFOJq8nqrsa4kPhRRwSxkRxHLsU2KFGjuiy8qy4MTG7RIPuy3PgjhVuzT3RfnpcqJ4vgWI6EnJmHhKO413RfRKSiP37yJYyjtEc5SW4lZh4SiOPdF30SbxXS4FstieK+IFuXIlZh4ehDVcCd54jv2IS0qhvwYrpUjkijDjsVXAneUnSIqojyxrukQHyRRwc5Lokt8pcGF8JxlEjlZRKFWPeIzA3jTHcRHwT/nO2+BKjFhaKGYU/lkbxMSPzRIT1rKz4hbGLhat0NDRDEa2fBJWjDxNPtlm3QlfOWJhqZKGnZjVim1tIjLTuuCMtWbdCj3llKCnyTwnA2lsxSlhfwQxFPovshKt3k4qXI4OPBLDUhTlhPchiqXRzwJVm4WTwHzE9OZDaCJYlEsRy2RDBr4hRo4ys5KrnOWIokpyxHSFFR/kWG5byEkuMrHucc5zxEluSm8RnHBDDciMVHKyrOOcpz0jfzSHJzEhJvgw8PRlY0mcfFliT1e1EI7GLP5Vng4fzPNqxOtpEpaVZh/WzeQ6iiUtTERV7ZtCfZk92ojfZCj5ynvIgLkWVeC+wuC/GbyZhcZV3RFnEmc8ZzRHwSMKVMQ1XBL3ojK42c89GJGnnhT1KhquDVolaNSKvd9GNh3us8OejZ8E4d4mHi1tI1XwKPd9E4KfJPDcMk3DgTv3RIYifJd8CWnpxMC/hONmP2bow8e9makfFwLbjplBSJ4Y04PYhjCmmfEcdPJSFKoI92I6Rh4Kjz+Q2ok8TYb1PchC+CMFHK+j+STcXUTExNJep75YeF3ZVdCOSc9MtMST0byHLW7eUVbIYaj0I/knie7TFkMNcmLiqGxZZhR1Ppe63NWqVdiMcsfE+UsizBjtfQ6rcwd7kJVk3Sssi9jDfQ1a3FL2HCzxHRqtjZhPd5RJKz4nb6JcF+8kWYctUcmlyL2YldOJHUh7ZRm4uyMlJWYkVyYM9MqfVjYdbo3LZhY1bMxElujBxtLp9TVmJhuHA2xNp2hXOJh4rw3pkX1TgpGJCcMo8bkJF9eJha0PBlBlUhTaFO+uOHqiiMVHjrtIczcmtWyMP8Ax0t5HHW2X4MT3EYNvYw8JR68TEb9sCMFDfuYr1MohHUQgodWNifLEwsK2TksNUPd2xEIamRioql040/lRDCpUInLSrG7d5RV7HHRiOokY6Y0IfBiv2iHwQXTxFDzlnD4sojH04ifI90Oz/HlvWTMWNqyEtSvpxYFDMGel0zkxMPwYU72fVi4dboZRhTr2yJ4XgwpuPtl1cmLgd4mkjKhpYi3IuWHt2FJPjqavkxP8fvE+HkTEy+t7ksJdine5/ApUJ304fwrpe2TnXA/vlo8kYqPBfVriNjkOVkcNvcjFR468bES2FpitiU7yjHVwYaUV9+rExNOyIxPVjWxKWp3nh+znpb0qyFyetl0a0uTGlqdZRMOVt0J30P3TSGcGva2Tnr4Ip/cl4NWnZl+c+w8+eBzTelFMofseoUtatEcpcdDfZEkR4olEj7XZHGjPYWzp5Q9ktPQ34J+2I0UULH0qi7JJwdojLUr6X+Jt2MTC0ZrF0rctYv8mHiadpdTd7IngprYktLpkXQppr3CxKZCamrXU3R6ae8ieE47oU/ImnwTxtDohirh9V0KOv3SJRvglHTyVRLElFbCxt7IzUsofCuiU1EeJ/8ApBPuWhRchRUTnZnGz6bSMTG1bIjFv3SHOuDeRDC7vJrTx1YuNp2RGPeQ5XlGLkyMdKGrE+z6Jy0oXJiSr2xEqzwod3l8H8dGI9T0m0R/VIdzdvKh7KjCjpQ13QneeGuZZVq3Z/kb0ivsRX2HvKhRV8Zfzl2JcjOeDhbCir4Kymv4MDZDWndCdnKzb7C2JJHEia/jJow36kdxOtmYi+ZEXavJuhI5JKnQ88GS+BjXZifpsWfxfwcDV8k4aHnVboUvU/kw8Ts+i72RxxlOGpEouDE6HWJyKUsNkMRS6G6Ixrd5zwtXB7oOmXGSpmJhuG6MLG7Cknm3Qlq3fQ4WNXsTwu6ITcXuayHwLJtIlMbc2Rioci3ftIw89HJ8ObnRiYl7IhDTvIc/BGLkQhpzsarjoxcatkQj80htvKMdRGOlZtaheHlJ6Tl2TejZclFFEIamLbbP4f4ynLSiK0q2JXuzGlexRX2FH7EI655tdxOzEex8MaF7t3libyEiMf4FuxLKrPh2eT5L1bISoZ37H/4Mn/Rgc5NVuiLvJvshKs5fyN7Df3P7MGVOiSsT+VmG9L0sboWeJHUiy/uf2X9yElNUT22Zhzr2vKtX8dEo6kSWl1Z/Z/Y/KE9a25IYnZ5c7IW3HRJalRODgXQ6nyJvDZDFvJuhRrd9LWonhuHApeScWnaIYlimWhLVuy+l7mjTuYmFq3RpYq0xHLwOVEpa2QSivuKDfIlXVzsfDsSmTn2IRXMhyshh6hKulDi1vEUjFxSPudseUIamRjpXRY1qHJw2ZJuT4G1hr7n8lFfYUb7EIKK6XcN0P3vU0Rjbtk5aUclfYr7EvajBjpV9DjZvOW6N5y34yk6WSRwuxDjsRyic7MWpOuxNtypCVZSO/Y//AAsk/ujBfuHk007iTnToiq6Jbd0RkN/cv7l13Iy1KycbHdaiG/ufTiLS7G67l/cv7kZ6XybTRpkmYc/U26px1Il7XVl/cv7l6XaIv1OOT1NO1kaS26mrMTD072X9yTTW5GWlkJka5L654V7j22kd9jDbaExTv8hxUj0kJ+1HJiGFhyk7Qo1+Q5UOVkuMo2yGF3f5DlpG9RifERs3IQcmRWnqtJWYmI8SQnpjqZKTk7NyijCw63fV/kT20oh7VQuDGlqdFfY0vwKH2FHXOhdHBh95kcsfijSKDJR0ojhuiKpZLKXukjiWbNG/Y0fwUSj/AAYW0s2/BiRaqSE76JoW0iUfuf3lgS+UZL6WYUvlfTKOpFdj+z+z+zBxNLpmJdWi3F6kRlrVrqxIah7dzbyMwtpE4rFWxhYjg9Mi+vEwu9ksouNC2FK/yJQU1uYuA48GE0uS7e2SlQn+RDhWK+wofV+S55WvI5/cjDU9jDw9C66G6G/JKSXDHucEI6+4lXXiT9R6UQw+7MSWsrLYw4Xv1N0rIrU9TIR0oxJaFtl/Ql9h1FGBGlfQjFewo0lHJGNu+BR+xGP+pNdkjT/rmuMorc75vkUf9Sv9Rr7Di/pIqpcZPKSuIsnk9yaa3oab7FMpkW4sW+5NWS2lqF04q7js3Hlhz1LSzRpZF6Hvwc9WJC90O/JX3Ft3IzfklFT45Iy07SYuvFwtW6KruKTj3FJPmR/Apfkzwr3RbWzYnFdz7osUuvDjqihJLjr/AILrkcryft4LbI4bumJV13Q3Rfkcmu5bfc/sUJPdEarbrxH2IR8mJiXsmX9z+z+yKvhkHarqxJanpRHwizEkpM2FXkVeWS90qE62fS/dOjuSdDaXxEqchafuR0/cfxHt+5dxtdG95t6TVpVyKi+xS+kaVcDS+kpJ/CRmpbIi99LyXBHjJ5XtZSa2iLdcDj/qOP8AqafsRxdCpmremONqiD236LoSvkXhocX4Kfgp+BWt0j1I1uTjZhyfD6pP5UYmDXBT8FPwbkJSMRqKt8mHLVt1ylSPS2vuSjKPIrQpSY0a9K3Fi6laE1Lddajr9z4J4b+UuXdmxwKVEcbXsQn8r6Iqop9XBKWp0h4jbqBdlPklK+wo32IYaQ1qE+qc1hqy5YjEthyfg38FPwQg3yhbcD9rvqbUFZKde5kZS5Nzc3EpMiqJLuhO10SdI+Hk1LCjcuTU5u7N/Jv5FfkbcVyYULeoasT7PKsod2XSF9bHL1HbZf8AsRf+xf8AsRe79w6kqcjDioxpD9j+2azXvdmOk+RaV8xa+obVcja+oen6iPtktJNXuiL1ETiTz+J0h8HtW1kaToenyx6fJ7R6TD/Eh/AnY6jK+j4nlixr3D0vc9p7TYaXYw8T5ZjVckJ6l0N0RVbvLEw0t6NvBt4NvAtMuxTw3Zh4nqLputyKv3PKUVPknDS+Cv8AUjKvlPj7E4OD1IhiUxSvp+N12zlCMjTp+UTcuw40Th3Rq1fyQmKV5YfwIfs/joboxJ0XftRGNcFx7ja8kIaiMdOcl3Rd9Ep0SbxJUJLDJSj2NjYhBSKrP4dui6J4tuz4nbNvBS8FLwUvBhwXNZv279Evc90R39zJN4ktRX2K+xX+ol/qT3dRRFUspx7ojvlN7bHCo+NmL8OxT8FPwRUvpHfeJBS8Hu8CGr5IunpeSyfuekW2xiX2Fr+x7/sPVR7/ALD1/Y9wuCXtepCJfFlJ/KhLTtk9XYnq5bPd2Y9Xk93k93kw5NPdk1W6H7lsQdrKT7ISpUcZbxdDvyb+Tfyf2NX3MOWtV3E6d2J3xnHf3PoxIOO9n/Y/7F/7G017pCbw5bEJKavoS1v7Dzasnh6e5a8il/sKcK5MWGndGFO9hSzbv2oSUVS6ZYVbpkZRXctSexiwrdEJ6WJlsw/gRyLb25OQ3RJ6mYcBuUT3Mhhv5upqt1nKXgxJ9jCjUbHKXk38m/kjCXS1aE+zzxsXshKz+z+z+z/sQi3vfT8DrLEl8tnPsMaVLQKvJt5NvItP1GyVpmElJ3eSyl7XqQne6NpTok7elCVGPJcM9nkWjyL0/JLTWzI+nXJ7M5R1IhLUR4JSoitOWLXc/D8H4fg9ung9n0j0fSe3wQ+EZH2vST7Mbrciu7zml3Q9P0iprdDUfpNvpNvpP+pF6oj9khe2Ww3SsgvmeTLJxtWcrg/6n/U/6n9G6dpDqa1ohPsll8b+3S1fJONPZG/g38G67Ek8RcGHNwYpa1ly9KONurEg/lR7vAnJdh6pqmSTw5EJWKQ3tsQWldco2fiIVv4jFhoZCfYsh8KykxuxsnKzDSu2SlESUiOGo9aK0kpE50QVu2Nx7I9vg28EIKXYSrpRNd0RkpGLiUcs/o/o/o/oir+USrjoQ1q2FPT7WN290L8OO57n2N/B7vB7vAlLwSbexBUt8lm36T+wpNJyZhqt3lPU2e4WsXqEnO6PxPsLX36J7e5Cl7NRh7+554l9ha/Itfk9/k9/kev6hqXkw+Mpq0W5YZC5+59D42Pd9QrUqsal9Q0/qN/qN/qMJ9mySsqXBF630cZT9jPvqP8Asf8AY/7H9kJ+nL7Eov5eDX8lkdlS6pK0Shp5Zt5NvJsu5OuxhYlbDltsYa0ofXPCXJ7fJcfJiaGtuSMqExMUr/IaUuSWEluS0VlqIfAhyzlxkpuqIRkxKvyLocrylyQk1wWy5GHGT5/Ise3BiciLfk38m/kVvuQjS36rJz1z2FUtjHxLelF/c/s/s/sW29mGtcurHn8pq0wSZF2TemJt5Pb5Fp8ns+olVnt8mElfRiSqItXpEJWs8eu4lEqAlGmVDwyo+D2+DAarbKT8GHc4tGC62E+iUVfBTUuCUY+Cl4NvBt4E6d0Xas1NOmL2TEy8mrylHWqI+GV/qf8AUf8ABT8ZYEm/azGjTtGFialT65RUhpr5Sn4Gn4GYabkVp3P4L/InC1sOMl2JJiIwlW+alf5OJhKZPDlHkoi/as7S5J6X3KIYPd/kt0N3lqjVDoWk9pDDi9zjqvJ7GrTyYlN7LL2+D2+DbwQjGrrp4LMV0RjSP/XD75L+C/8AUv8A1E/9TEfZIwlUeMkPPTrxD4sQpMxnWyLl4Ll4Iuf0mqXeJHVq2Rc/pE33XRPdbErWGQ4Kynq+UXqn4wtfc/FH6o/UMPVe5WWDs2hLTN5VlY9fyk1itEHKth+oP1D3j1GA9qZiK0SVqyLtdFZYkWvci5S4Z7/J7vI9Xkow9SezHHUtzQ4yEX1SWpbDjJdxqXkaI2ndlOXMhOtjn8mcNZOGl02KK8kf/wCiopc5qX5MkpbM9GJH4UcjdcI1fY3l2I4aX5LlRYlZqkuw5t9jfwb+DDi+6/I5OCn2HKaPcypHuKmQU+/5GmTdsUVL3GI5SZpYlISn5FGfk98eWRi5ytZV0SexhR0xtkV3yxPdLZlP6hRf1CjL6imvmIRfOop/WRX3voZNe2hbLPESfLo0x+s0x+sSje0iofUNQ+ocYfUYelPZ5x2kT2n0zSfJWF9RDTxY1h/UNYfkejyPSYbjF2PJVB6elnKplaXpY1ho/DHoPaewhLDRKKxFZFxg6F1zw4y3HoPYewTgKWEuBPuhb/kyhGXJOMYOqPb4FKH0nqR7IrvknRs/yYL2qx6ux7vJGEmJafyXLJEr7M38lPyaX5IYb5v8njcvySr6j+yl5Kj5FGPkUIvuJUq65OMtmxLQqRiOK9p7PJUPJUPIlh+TTheTEqOyMKMUtS6puPwsaqOkTG6VlwZ+GfhC9Efppe0j6NF4PgWlLboddyfAsr3oxHHurNUPpNUPpIuLeyNUPpNUPpHKP0kZK/hHJVeXcxezFm3pVl2tzWvpHL3fCOSXyjl/qOX+pf8AqX/qRlcbZe1k+NRF2ujnLE3jqFLbgt/SW/pLfgt+BSkuxGcn2JKtxe5bdd1uS+HVRqf0mp/SW/ApyXY9ScvlKo5yi9Svrf3GpNWj8QUsRCliMcds075E090JqStdS00rYop7WQwkuRbbdcpKCHiOMdz1NSy2jyScGew9glFkMNR3PhddcmoK2PFfYttWyWJBjcS4lx8Fx8CcPBGMaI7e0fTJ6dxaZ70PGeq4jnq3oteC14NS+kUl9Jqj9Jdy4MNbbkdnpfTH3S4JO2J8zYpzuzU/pFJ/San9Ipy+knJ+BTl9Jrn9Jhxe+ojs9DzV6tieTdbkVs5Mw1iR4LxfBeL4E8S/cjVi+C8XwXi+CTxfBgpq4yI7e3KduGwuM375aTFg5rYisVKiaxWi517R+sP1T8Q/EJqb5MCd+1kdriyOq9+mXuelEo2qKlBjWI+GVieSsTyVPyVPyR9RdzFU17myGJvqPv1P3PSMlGXyn4hWIaZi9RdxKb5Y1XBGbhKpF+nK+xzv1P3PTlOGruPDku5T+oSb+YpZPdUQk8KVF6JbCkmPow4qS4IxUeMmrL6bok7Yve7yft3HiLujV9i/sX9iMUsmtSE76eNzEncjDhqdsc3HsObfYuXguXguXgTn4IX3RZLdWjlWLocpp8GLKlpIqUexcy5+C5+Bep4E8XwYk5NUzCWJHfKavdClqV5v7ENVe4k72MX4dKEpo/EF6p+MfjHvctisXyVi+RX3MRbWhO98o/ETyfudHY0Yn1GjE+o0Yn1Gmae7NE/qNGJ9R6eJ9Q4T+ow4tStsxF3Rdi3iR2WUpaVZhqlvl6cvqHhSfzEE1tZ6UvqHhP6jR/saP9jR9xrQ7RLdLEJLX7kxZuWlWYard5YsNW4vcqscK+Y0ryaV9RpXk0ryKMXs2SXpujBna09LdKyKqN5vDfk0PyaPuaPuKP8AsRil3MSGrdGG79sjDmc9DdIitKHlKCnySw4R5KwyPpGqFclE46kJ2tLIStCkVnD4FmmPZ50Nk5UjkiuyHceBzl4Lke49xFVz0S9rvpxJ0iKc3Q4yj8I3M957z3lYhFT75o+B/bOySfyltK5FOb1FT8mmfkqfk0z8ihieSsSO7ZTxJEYyjs3m/ZLOScuCXtiQXzGIrlyaX5ND8ig/qPTl9Rokt9QoOTuz039R6b+oWXwSrKK9xPkb0ogqQ+BYcPqPTh9R6cPqNEU/iHhxb3Z6cPqPTh9Q8OHkjGKfIxe10QEqdZfHKvGcoYd7mjC8iUIy2Y4YfdjhheTTheSsPyVhlYZgNbwF3gyOmPtWb98qz5JxUGVhtWz8I/CPwz8I/DPwmiMtLE9XR/7JfZDHk1ezHhRRph5NOGVhi9ITw48GLH5kRlTIs5yRH3yvsPocVLknGMexcPAp4fg9WBV7mLGt0QlTExM5yg/aujlEZX7Xk5Fk5WzCiNNL2jcz3FSFGTIRrnpe5B17HnJk5amYcPbY1LyaX5NL8ml+TQ/IsN+TjbJZSWpEHezz0O+TGlb0I0fc0fc0fc0fc9P7iwl9RNaNrMPCT3sSpZtalRB9nlGKctRP3yo4Q4xfc0R8miHkWHh+T08PyOEY7pkYYb3bNGF5NGH2znHUiDtEK1E+T45ZPgXon4B+AL0b2JelfuPwD8Afon4R2JqzCdkqUyUqRBaVnPTzI1YJKWD2Lw2rY5YJeEasMvDNWGa4p3EnvTiNxS1idkpaUQWldE4pojJcMcoLsa4eDXDwa4eDXDwKcPBiVJ3EwZ9jnKcqVIgtKrPjJpS5JRhHk/DPwy8MjPDQ8TDcaGqZhy7CdC3MR/IiKUVQ+qft7Gv7CxfsLG+w464klpdGHK8rNTIfCul1djeU5URWp0NbUh6vJT8ml+RQb7kI6evEj8yIvUrJMxJUQWpjhXc0/c0fc0fc0LyLDT7igoZLfomqetClfBJRl3H+HGyKT5NMTRHyaIeTRDyaMPyenh9h1KW5HDhzHpn7XqRqVbi04cbRBdzEaS3PwysMrCEsErAJenHgXoH4AvTfw9GJ7HqRhU9zFe9IiqVZPjcU8Lwa8Hwepg+D1MK+CUsNP3HqYPg9TB8DnheDXh+BO42sk9EzFpUz45dDPVh4HiQ8EJxfY9WHgeLHwepHwepHwepHwa4+DClqjQva6ZGduhe+Vl9OKtIpquD1Psep9j1Psep9jX9h4lqqPhZhytDIe+WrraUuSThE1wNUDXDwLFguxjSU/hE6IyssVN3m11Tvsa5eD1JeD1Z+DFTl7qIumJ5w+FdF0Xk2SdmHGzT9zT9zT9xYdkI6fyW/A3RJ2yEU1uaYmiJpiaIGiAsOK3OSjjpvTPSLDj8SMWetiUKKgaYFYYlhiWCYmmPwmGsN/EJJcdPJGtWlk1TXgRiyjdMvDLwxPCFLBNWATcE/sLEwT1MEi4S3j0S3W5/jdzmbbzeyFjQ8Hrw8H/kQ8Dx4eD1Yx5R6+H4PXw/A8eHg9WHghJSW2U1aon/6jCaSLRZZY8ZR2o/8iPgeIpS4PW09j1/set9j1vser9j1PsQxfeShe5jPStjCa07Z2Xk90W4yHi12PVfg9V+D1X4PUfg9V+CT1OzClWx8SoW2xfQ1ZpOCkxzgux6kPB6kfB6sfB60aqssK8rE7zfTZJbbDlNdj1JrsTxW1Tyw+M4/CLN5yyh0YX5Cznx+QvhELqn8Qv8A1/kTI89a/wDYT4I8GL8XQsp9hZYXHRIwO5L4iIiXHS+enD4yRifAQyQsnlPnr+Yl8JifAYXQs8Xkjx0vKHIh9bFyT5yWUssHvnEf5Mxjyws//8QATxAAAQMBBAUJBQUGAwUIAwEBAQACAxEEEiExEyIyQVEQIzNCUmFxgZEUIDRioQVTcpKxJIKiwdHhNUNwMFBjc5MVQERgg7Li8SVk8FSj/9oACAEBAAY/Ana5z4rbPqtt3qtt3qtt3qtt3qtt3qtt3qtt3qtt3qtt3qtt3qtt3qtt3qukd6rbd6rbd6rbd6rbd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6V3qukd6rpHeq6R3quld6rpXeq6R3quld6rpHeq6R3quld6rpHeq6V3qukd6rpHeq6V3quld6rpXeq6V/qulf6rpXeq6V3qulf6rpX+q6V/qulf6rpX+q6V/qulf6rpX+q6V/qulf6rpX+q6V/qulf6rpX+q6V/qulf6rpX+q6V/qulf6rpXeq6V/quld6rpXeq6V3quld6rpXeq6V3quld6rpXeq6R3quld6rpXeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq6R3qukd6rpHeq23eq23eq23eq23eq6R3qtt3qtt3qtt3qtt3qtt3qtt3qtop3j/AKQu8f8ASF3j/pC7x/0hd4/6Qu8f9IXeP+kLvH/SF3j/AKQu8f8ASF3j/pC7x/0hd4/6Qu8f9IXeP+kLvH/SF3j/AKQu8f8ASF3j/pC7x/0hd4/6Qu8f9IXeP+kLvH/SF3j/AKQu8f8ASF3j/pC7x/0hd4/6Qu8f/JW0FnVUDVQAIayGO9YOK4rKqyK2lmP/ACY7x/8AImLgs6rVaSsAKrF1FUk0VB6rDkvcV4BDx5bu7cqjLeqg4rgViSO9YOqFuKoWreFg4f8AkZ3j/v7FwC2r3gsGnzWq0LF1PBZnzXErFYYDiu9Vd6K63zK7lePkg3jyPPfTlcOOK7xyfL+i71Q5rDEcFUKjh5rDFcCv6LVeVjRYsr4FUIIW2sCD/v8Ad4/74xcAtqvgsGHzWq0LWkp4LNzvEqpWqFiargF3rHAKg9FreioMSq5lXW+ZVAqdVvIX+Q5AeOKd4cjXcDyV6ruS6ctxX81ddn+qqMCqHArV9FQ5rDFcCu0FhgViKrA+S2fRaryPNbVfJZNKxYQsTd8Vg8f75d4/7yxeB5rar4LVjJWAa3xXSflC1nHzKwxXBdorguJXZWOa4BVPqVhgOKr9StXLjyUZ+ZYK4zPeeCoFcbtH6KgVBtOwCATkAneCb4IjihXPIogotO01UKuO2v1VCrr/ACcsVrYt7XJ2m/VcV2hyYG8qHArA18VrYLA18VrBarlrNWBqsKj8JWEp811XLWjosbzfJYSBYH/eTvH/AHZrPaPNbd7wWrE4+KwY1visZg3wCxc9/iVU0CwF5cFjiVgKeK1itVq1j6KjR6LE08OTshV38StTHvVTrFUzPAKr/wAq4Lsx/qqBXGZ7zwVAqlXnbbs+RztzdUckbeLuQpnhySM46w5BKN2DvDk4OGRVDg9uYVDiFR+LNzuSrMuysPRVabrlR+HfuXfxWOuO7NcVqmvcVRwu+K1TRazfMKo+i7SxFD3rA+q1mrVcsReXZK3FZFvgtWVy2g7xC1ox6rFjgtunisHA/wC7HeP+5tZ7R5rbveAWrE8+KwY1visZg38IWL5H+ayAXFYCixctVtVwWtj4rVb6rElUAx7l2VU58StUV71rHyC4LK6FXM8SqAXnLX9FwC1MG9pd/FYqr/y8mjj2t54Kg5NIdgbP9eTDaOA8UG8g+VvK3kik77p8+Uwndi3w5L7MJB9VUeY4KhxC7UX/ALVgqjVfxCuyYO47iqHFamI7JXA8Cq5HiFrC8OIW4hahp3Fa4u9+5V+oXaCocPFapurEV8FuqsD6rWatU08FuK1hRarliKrsrOvisWei1ZHN81hLXxWLWuWtGfJYkt8QsJG+qwP+5XeP+4NZ4Hmtu94LUhe5YRtb4rpafhC1nPd4lYrDFZUWLlgKrgtYrVbXwXBY/VararE08OTVb5laxquC1W0HErW1lisrg+qrSp4rv4Ba2qOAWAoqUvO4BVk/Lu5LrRefwV52s/jyaOPa3nsqg9eTRN2Btn+XKT1IsPPlmf8ANTl8z+vI5vEJruQPZ0jMQg5pwPJpmfvN4oOaag8lW60W9vBAg1HiqHELE34/qFUGo8VjnxqtfXb2gqgg+aqDddxBXOCo7TVgQR4rVN0rXH7wWYcFqOp3LWHmFuK1XeRWsPMKuBWDvVazaLD6LB1fFazVgfRZ18VrNWqaeCzqtZv0WBWQPksnN8FqTuHcVm1/iFrQ18Frse3yXSAeK1Xg+f8A393j/wB61pGjzW3e8FqRuctWNo81i4MHctaVzv3lur4rBv1WYHgsSD5rVaswPBYkeZWqFmB4LEjzK1RVYuA8FjTzWrrLFwb4Ld5rV1j3LEhvgt1e9UzPALcwfVbq8SsSK8FuYPqt1eK1iAsNRvEjFYZ8VUkBamq3tELD15LsVKb30WHqv7LRRbe802VQetM1/ZBjMZX5YfVBox4mma/si7M5AU3oNzO803r+yJ/kmE5u1sl/Zf2T+553L+y/spou++MOK/sv7K7/AJcuI7jy38dC7a+Xv5N6vxAlvWj/AKK801C3q/DnvZuKpi14zaVvV6MljvoVdkBjf9Ct6q0lju5c4D+IZKoNQqirTxC1gXji1YGqriDxC7Y+qpiDwK7+IWBveK1qt8VX61WBr3FazSFx81quPmsWehXesHEeaxFfArWFPFapp5rcfNazVqn0KzBWLfqsaeq1aLVkePBy6UH8QWLGP8CteJw8FtU8QsJG+qwP/eHeP/dNZ7R5rbr4LUjc5asbW+JWMwb+ELXnc9bI81mB4BYkLVCzAWLq+K1cfALcFi6q3eiwHqsX+izAWrj5LF9PAL+qwNT3BdgLE3vFYuWqKd5Ws4uXBalXLXf5NWGCxOPBb42/VYVrxWJXN1p2jkrxJc7iVvV0Vc/shXpST8u4Leqk0C6zIfq5UFQFvWhiqZN57KoK954rei91aBGaQHSO3dkcFvW9BuNyHE/iW9b0+lau1R5oDHBb1vU4x6Qret6hkxodQret6LcQcweBWIo4YOHet6oRUIRmuidsHh3culhGO9tdpVHmOCy+qri1wycCrkwpwfuKyVHNqFqDSM7JOIWHpwWSvR6h4blSVtzv3cmzjxCy0g+qwz4FYtBWofJy5xl3v3LcQtXUPctkPHcqYA8CtkLCh8VrMu966rlqm6sWtd4KhoPFYUHgsCD4rWbRdVYOWTT4LWoPELA08FmD4rFvoswCsHrJpWLaeS1JKeBWE9fFdRy1ofQrEOb5LpB5rB4Pn/3J3j/ttZ7R5rpK+C5uJ7lqxNb4lYytb4LXnc7zW7zWFPILADzW2B4LFw81q4rMBYvqtoLD6rGQDwWJHmsDXwWYb4rF9VtALVxWMlPBZ4962vRYavitZ95Z0Wrr+C1n3fBYZ8Vi+i1PUrXeXfos1i7HgFno2/VYHHis1djq936Ksr73y7lmql1Aubq1nbI/RYVrvPFZlYk9w4q/NlujW9ZlaKGpl+jVQEknEuO9b1mVex9nYcPmK3renPNcFrV0jtZ3it63qzR44vvei3ret6tQx2h+i3rrJ4AdezHimPFdYLet6E9Do36r/wCRW9ZFFrgSCtBLUnqO7QWRWS0sWrJ9HeKIulsjdph3LJULahaoMkXZ3hXm4hZKtC1/aGa55t5n3jf5qoFR4qhaqxavy7ldlZozx3FbKxZ5rV1xwcrpbcfwctlYC4e5YsEg7s1hnwKxYCtXDuK1o8OLVhQrZA8FhQ+K1o6d6yaVgLvguq7xWuy4q0aVgaLZa7wWsLvisAPJYO9ViwHwVDQeKwNPBYEHxWLPRbq96wNF1SsWrMLILADyWrK9v1WErX+K14mu8FrxOatunitV7T5/7R3j/sNaRo81t3vBakL3rVhDfxFYyBg7lrSyP810X5itlo8Fj9SsG+i2APFY/RYgeawbXwWyB4rE+iyAWAqsg1Y4rJoWqyq6rfBY63isaBarKrFwHgshXisaLVZ5la7q9wWAAWJCwaGji5a5vrcsSFgAwcSqnWdxPJSuPAL7pv1WGfHkpm7shc4643sNVG0AWYV0a8nZCvTkH5Nw5M1cZrynqrSSOvynfw8Fms1ooqGU/wAPeqB1XHEuO9ZrNCyxuoXYvd2WoNbg0LaW0o4b2qznH/yW0tsLaWfRx/qf7LNbS2laRe3NK2ltLaU9nLtl15vgVtLaTmOdVpFE6zyP149/ELaW0rpdjmHDcjFKaTN+vetpbSD2vuStyctHJqTDdx8FtLaWkifck+h8VcfzcvDj4LaWavQPufL1Srj6xycDvWaxxXMvp8jsldkrG7vy5KOFQubeadl6pIDGe/Lk1hVajy4dl65wOj/TkxBrxWq68ODlrtczv3KoxVaEHiFgb34lrsc3vzWGKyIPcsDe/EFrxuHeMVhisAW+Cwx8VrRnyxXFYAt8Fhj4hYxnyVKeqwBHgsMfELGP0WI9QsBTwXHxCxj9Fi2niFgPRcfELoh5LFhC1HuHgVqyk+K1o2uWvA7yWteZ4hYSt81g4H3XePJrSNHmtu94Lm4nOWqxjPFY2i7+Fa8zneaqXfVatVnTzWLysT6lYEnwXDxKxkPks/UrAk+Cww8SsX+nJteiwFPErGT05Npao9VrSenJi5aoPiVrP9FXesTRagLlrOp3NWGfJqAvPctd10cGrAefJQVc7gFjqDgM1gPPkxxdwCx5pv1WA8+SrjQLAGKPicytVuPHfyVOAVIRcj+8I/RarfEnMrJZIxWcY9Z+5qwBJObjmVkskIom3pnZDh3rIuedpx3rZWSrdq44NbxKq8XpX4vK2VknOcKAYp07m60xveW5bK2PoslapKde76LZWytlSaucY/VZLJZKzzU1X807+SyWytlNtMbdePMcW70HtxBWSyQczVlZi1yNW3ZG4ObwWSyQwuuGy4ZhaGcUl3Hc5ZclHN8+CpNrx7pf6qoxCyVHMqFhz0fDrBaqyVHNBC5o1b2HK64aN/ZdyUIBVYXXPlOIVJWXPmzCqKELcqxnRnuyWuy98zFg4OW5VbqH5V1ZB6FUOoeDluVaUPELBweODlrsLe/MLAgrEBar/Jy1mflWYqsaFar6fVZB3gsdXxC3FYOu+CzDlrNIW0CsMPBYPr4hYivgsTTxC/osJD5rc5YgjyWYWDyFtArELE+o5MHkLUtDvNbTX+IWvCD4LoCpm6YtaHkaoWvLI5ZLZWSwjKyosbxWzRYNJ8lsXfFY18lsLInwWEfqsfotknxWIotWNxWV1Ygu8Vs0WALvBYMu+K1qlYMosVqxHzwWsfJq2FktVhf4LHUHctm8eJK2VjnwWEdwcXLXq8962ViFSNl/v3LnD+61UDaLJUzd2RmsRoW/VarfNZKpwCpAyo+8dkrzuck4lZLJXbt55yaFenpTdGMlkslU0A41VGc3Z+3vd4INY0ABZBbkI42h8zsm8O9Emj5HbT+KyC3Ik0AC9qeNUYRN/mty3Lco7IP8zF/4VTBbluRcaYJjt76v9VuW5blH80R/VblmFmFI0HWzb4qOSo1hwWY9FmFn9EYCeak1o/HeFms1n9Fp4Tzzf4hwV8HxHBZrNXX/AP0hHO6oOzLx8Vms1iVes51d8Ry8lg6jhm0jELNbSvXrknaaqWjZ+8aMPNVD6hbSo7WC5p+kb2H/ANVdJLJOw7NZlZq9G4xu7svRc428O0z+iqyS8s1jnxWq++ODlSS9EfmW0VQ4rm3uZ+i1heHFq28eBzWZVcjxC1ZL3c5c41ze/MLVfXzWOK1Xub5rtjuNFrEsPzLNcD3FYSV/EtZp/dK2vJY4rVe5vmtzvotYFqwcD5rh4FYSeqxFfArHV8VuKwcR5raDli30WJHmsMPArB/quqfNYiizHJLhXWOSwZ6lY4eCxx8SsgFqsJWyAsSVshblhH6rcPBYi94lZALDW8FgwN8StY+iwaFjT1Wq28tzVjreKyCxotVlBxctd/k3BYNC3Kg1j3Lqx/Va2ue9bljRc22/37lrvoODVqgBblrEBajbo7TlWR2kPfkty3Klau7IWJETeAzWqB48mYVyHnXcdwV6d+kPZ6oW7kqXABUh1GfeEfosMSc3HMrNZqr3eA3lB9o1Wbov6rNZrNCKLXndu4d5RJdfkdtPO9ZrNZowg/s8fSHieCzWazRJdQBSWt2cuz+Hcs1tLaUlHGrtUeaYwHACi2itorNWQ13OCzWZWZWatFnrsPqPAraK2isyiGmkjdZh4FB2TsnDgVmVms0bTFUt/wA1g396D2uq05FZlZlFrsQdyuyFzrP1ZOz4rM+qzK3q8HFkoyeEI7RqP3O6rlmeW9Z33PkrqlaOSsUvZJz8Fn9VmqPF5ajtMzsuOPqruLX9l2fLXZf2mmhWI07OIzWqceBz5MRVc07R/oucjvDtM/otVwPJi0Fc2/ydiucjp3txCq0grcq0APEYLVcHjg9c5Hc78wqtLT4LctXUPyrNknjgucbc/RapafBYhpWo66uq/wCi1hc8Vg4FYhq1ZKeOKya7wWtq+KwLStwPctWT1WIB8CsdXxWYKw1fBYP/ADLFoPgsdXxC3FZKXLaKwZVZNasTVbIW5arKrqhY63iVgGhYkLVZ6raA8FjreK3LMLVZ6rF1PBZCvetyxIWq0DvcteSvcMFgAFuW0K8AtUBo4uWu+/8AoqCgHgswqVq7gAt0Y781Vxvn5uTNUvXndloxW1oh6lVzd2jms1mrt68/stC136JvBua1cFms1cBvydlqrO+jfu2/zQDdUcAFtLaVxp0kpyYEH2h947mDZC2ltLaQjj5yY5NH81pZX6SbjuHgtpbS2kIojfndkOHeUSXl0jtp/FbRW0VtFNghdz8n8I4oRsJoFtFbRW0VFZWuNZTrfh3oNBIAW0VtFbRVjhqcX3j5LMrMrMrMqwmu8j6LMrMrMrMqCWpuyjRn+SzK3rfyCXHQzYO7ncfd/wD1Xn8h/ot/LdOI71vfZfrH/ZAg1B5S17bw4LfNZ/4m/wBUHMN5p38myqPYCFgNPFw6w/qrzCDy0c0HvWHPx8OstXMZg5hZLJazceIzWFJ2cDg5Xdl/YdgVlyVLRXiM1qkSt4OzV140TuD+WtKHiMFquEg4OVJWmLxyWFFuVaUPEYLVeHjg9c4ws78wqtc13gtyrQA8RgtWUHueucZTvbitVwK3KuAPELVkr3OWszzbitoV4Hk3DwWrJ+ZYtB/CVQm6e9Zhbge5asvrisQHeBWtq+KwcCty2j6qWjRtFY0HmtVhKya1a1XeawaAsaBarb3gtkNWsb3msGgLILAXvBbAb4lazr30WDQFkFuqtWMDvcVrur3DBarWhZBaxAWpHhxdgucf5NwWq1oW5YkBc2y93nALnJMOy3BarWhbluVIxpD3ZLnH3R2Wf1VGABbluV0a7+y0LXcIm9lufqqMACzCzC13juFMSs/Z4/4j/RUZQLMeizHoi5z2gDeVzR0UX3hGJ8Fq5nMnMrP6LNZoxWYg9qSmDVg6rjtPOZW19FtfRbSEUWvO7IcO8okuvyuxc871ms1mi9x8BxKdPMefkz7hwW0tpbSreUtrJwdqR/hW0tpbS2ijrdDH+q2itsraK2yrCbx6VbRW0VtFbRT7pN9mu3yUcgcaOFVmVtFZlPjeTRydDK46aLVPf3rMrMrMotdiDuQs8jiYXdE8/oszy7yr8VXWfrRjq94Qex15p31W/wBVv9Vv9UZLMbj97K6rkWmscozYSt/qv78l9pMUvbarlqbd4SA6p/ov7r+6/uqkEO3OacViPaWcRtKrDXu3jlo9gcuadpG9iT+quyN0L+DlkslQsDu4qsTjGeycQueiw7TMQqsuuHcsgtkKrOaPyrFjZh3YFUOo7suFFkFkFW4AeLcCtVweODx/Nc7EY++lQqtukdyyWLAVqSEdzsVrxXhxYqVAdwdhyYtBWoSxdWT6LXYWeIWqQVksNX8KweHfiC1o/wAuKzoeB5MlqyHzxW030U1S465WDPosiqYk9y1YyO8rWcf3QtknxWRWK1WOcuwsQ53itkrIqmJPALCO6OLlrlzlgyiyKqcFzcTnd5wC1yR3MWDMeK2SslQNL3cGrLRN9Sqlpe7i5bK2VV2A8VzMJ/E7AKs1ZO7cqBlFsrZVxrTJJ2WrnTo29hh/mqMjotlbKvOo0d5XMs0bPvH/AMgr1L8nbccVsrJZLRxs0svZBy8VpLTSR25vVCyWX1WSLnUa0byVq81ZuO96DGMDWjcsgsgsghDE0PndkOHeUSdeV2Lnnety3LciTQBe1PHMs6JvH5luW5bluTLOyl+c3fLemsaAGtFFuW5bluVsmw1pKei3Lcty3KynhMFmFmFmFmqVU1mr0L8PBZrNZrNMtjerhIKZtQcHAgra+i2votrBOjeagr2Wd3ODZd2wtpbS2lmjNZsWnbi4+CD2PqFtLaW0hUkOGy9uYQbajh1Zhl5qt5bRWaIOI71WzP1funZeXBXCTHL2HLaW0VtK+ateOu3ArXrPH2m7Q8lVkl4LaK2iqO1h3rmJXN+R2IVJw6L5uqqhxI8VgSt6vYsf2mmiz07fQq6SWP7LsFmVvVHC8O9c1I5nccQucjvDtRrVdjw5P7q9S67tNNFqv0g4PXOsdH35hVa68O48lHC94rUc5ngcFi0SDuNCqOqw/Ny1u0PELUk8n4rWhr3sVK3TwdhyYtBWrVngVgWu8VrxEeGK3+imDWl2uVuZ9VrEu8VhQcmLvJajPN2C1n+TVljxPLSt48BisGhg+Za7y9YADkzVIwZD3LWcIxwbmq7R4u5aucAubZh2nYBc7Je7hgFRtGhZrNazxXgM1q0hbxdmrxOkd2nFZrMLMK4znZOyxc9Jo2/dsP8ANUYA0dyzWazCLLONI7e7qhX536Z/0Hksws1mi57w0d65smCDtnad4K6zD+azWazVXHwAzKEtqwb1Yf6+6IohpLQ/JvDvKJc4yTO23kZ+5/Zexxk6MYzOH6INAoB3Lf6Lf6Lf6Lf6Ka1GtxnNx4eq3+i3+iyPosj6KR9DgK5KKoNXa2SyPosnei2Xei2XeiY6h1ZGn6rIrZPotk+i2StkqN9DdnbcPiFslbJWyVkUWltQU6xvBoNaI/KtkrZK2StkoZskbi143FGGVl20M2hx71slbJWytlaezCknWZuejRpDhg5pzC2VsrZRa6OrTuVYWmWDfETiPBXmCv8AJbK2FsKj4/A1xC12meLtDaCvMo4eKy+qy+q2VfaNHJ22lc9HpG/eM/mFeZRw7islkFshXoHaE8Or6Ln4sPvGYhXmFrh3FZBZBUexrh3rmZKDsvxC56K4O0MQqsLXDuK3LctdjT3rm5ajsyY/Vc9Ho/mGIVWOa4dy3Lcq0DXcW4LVe2QcHrnWGPvzCqxzSO5bljRap0Z+VYOZL44Fc60x95GCq17XDuWYWtQ+S1HmP8KweyTxFFzjSzyqFqvB8Fms1L+I8lBrHuWDAz8S13F30WqwBZLcqNF49ywaGeK16vWDQPBZLIKjRfPBq2WxD1Kq4aQ/MtkLJZBXWN0juDQta7C3gMSq3Lzu07ErJZLJXWjSP4NWuRE3ssz9VqMA79/JlyXGDSydli551xv3bP6q6xoaO73LjBpZew1VtJ1fum5eaoAAOA9zRRt003YG7xQltTtK/c3qt90RRt0s7smD+a0050k537m+HutjjGknfssRe83537T/AHQyMXp5MGNV2t55xe7ifdus6WQ3GJkTeqPdkAzfqpjeAp7sp4UKae73TIzbiOkHkmSNycK+6JYuniN5v9E2Ru/lx3cjZoTdtEeyePcq0uvbg5p3H3dNCdHON+53cUWOGjmbtMPu6WF2in47j4rRTjQzcNzvD3dJC7Qy8RkfEIMtTdEdzxsn3b8TtDJ2m7/FUtLNX71mSBa4OB4e5fYdDJ2mLnG6Znbjz9FVjweTPkvNOif2mGixuzt4jByoHXXdl2BWYWazCvDUf2mGhWD2TN78Crr+ad862gswswq7Lu000K1ZWyDg/P1XOtMXfmFqvafArMLaCrgHcW4Fak4d3SLnIyO9mK1ZG+CzWaqQK8Vzc58HYraj+qmwa1t871rC/wCJWDAFsj1WIHqtRt89yyZH51Wvr+JWDQFkFkFTBzuDcVqxsjHF5VZDpO4nBUDWBdVdVaxYPNakbQ3tOXPP0ndkFRrWtHcty3KpLQFSBml78gueeKdhuAVGhjR3LqrqrNquR0lk4NXPyBjfu4/6q6wNaO4LMLMLMLWcLxyaBiVrO9mj4DaKusutHgtpvotpvottvoi98rWtG8hEMdoYO3d1j4K7HQcTTEra+i2votr6La+iMNlIJG1KRg1Gkl57tp5GJW39Ft/Rbf0W39EGMdpJ37LKIyySX537TqfQLa+i2vottbadI+SjWo2yckSP2G9lq2itorbK2ytsp8l8mKz6rfxb1tFbRW0VtFbRVis946z7x8ltuW0VtFbRW0VaNY7KhN47AW0VtFbRWZRBJoVNZnPdegeW57ty2neq2neq2neq2neq2n+qpU+zT5Y5OWZ9VmfVZn1WZ9Vv9V7TZwb42mV2wmyMJIPet/qt/qt/qt/qrzSY5hsvC9ntA0c/jg7w9zJXXsqqSgy2fdJvb4oObRwO8LJZLZVHMBHAq9ZtZv3L/wCSINY5N8T1ksgtlbIV+Lmn9ww9FS1Qhv8AxGjV/sqtDSO5bIWyPRbI9FUso7tNwKwAtLPRyu7L+w4UK2QtlbKo+NrguZfh2JMVSeLRfNm31VW0I7lkFksWgqsJMJ+XL0WLGzt4swKu7L+y7Arcslkq3bru03BarxIODx/Nc9E6PvzCq0hw7uXXYCualc3udrBa8N8cY1S9dd2XYHkyUn4isTRc20v8Fi4RjuxVXVefm9zF2PBc3HdHakXPSl/cMAtVob4cuJVImmU/LkuceI+6NYNx4nP3Nd4C5qPRt7cn9FelcZnfNl6e7chBnk4NyHmv2iSjfu48vVXWNDR3e5fkeGN71zI0EX3jxifAKo1nnN7sSfd0UY003Ybu8UJbU7Sv3N6rfdLnEBo3lUYTDZO3vf4IMY0NaOHuhjBpJ37DAjLK7SWh+0/+Xvf/AKcB/O73nFuLzqtHemR9bNx4nkzWazWYTjUUhjp5lbQW0FtD1W2PVbbfVWgX27B3qCr27A3rpG+q6RvqulZ6rpG+q6VnqmvEjdHaGUOO8LpWeq6Vn5l0rPzLpWfmXTM/MnxGZldxvZFXZpGtlj1XYrpWHwcumZ+ZdOz8y6aP8y6Zn5lp4ZWvheecjB+oVfaI/wAy6eP8y6eP8y+Ij/MviI/zK6+dldzg7EIwWiVpplMMnBU9oZ6r4hnqunZ6rp4/VdPH6oyWSeOnWhLsD4cEHmUR8Q/Cip7RHX8S6ZnqumaqG0MB8VryNqMnDMINdL7TD22jWHitaaniFhOCuk+hW39CrmlF7hRXrNMYXdm6bp8kWTNcxw6wBLStaWni0qrJLw7mlZu/IVm78hRjcdI5vBpqFWB8k7Pu5GGvqgXRTMPAxlUeXMPAsIV5mkcOIYVsy/8ATK2ZP+mUTZnyRv36Nh/RAPhfK3tsjI+i2Jf+mVde5zXcCwqrWSkd0ZXRTf8ATKOls0rmjjEVesbrRTgYy5qpJY5h8zWGi+GtH/TVwtkDsqFqq2zTkfgXws/5FpH2W0R/O1lFes4ltDODmfzWvYp2O4Xaon2W0YfIrlJL3AtVRZ5iPwqj7JI4d7FeEdpiHc2oW278inP/AGgyJheaamS5m1md3afHgudt7Q7g2NVP2gP+mFdb9o6aTsRxVQLpBCz5miq+P/8A+QWv9p3B+CipZJgfnfFQIX7eL3dGqu+0aD/lhXIbe60S9mOIFVltAgHe0VX+IH/phX5/tM9zS0fogLPaXNj7crAPosftF1fwBXnfajmjiWBaOyW6W1S/LGKIG0WzRDgACV/iEn5Qrx+0JNIflBcUCLW+GHi9ovFf4hL6BXpPtKRo76LRWC0Tzv7RAoq2m3PB7LKK6+22gjxAQZ7dOHbo2Ur+ivyWqWzwbmOoXlfG2j1Cvy/aFoYO9wWi+z5rTJxc4qtot8pfwYcAmyPtM7ntyJdkrntlplmOUTDUlaS02uWNpyiBx8yvirR+ZX5rbM0cL2auWKSa4N7nfquetsz377poEbk87a4nXQiZPaZ7S7KNr0X2u1S3nZMa/ZXTz/8AUV+W0zjgNJiUW2aWVsfe7BqEc880/Gr10s//AFChBA+ee1uyYJDgh7XaZnynsvoAuln/AOqUZJJZu5ulOKc2KaRjOsb5owIOJldJSl/SGq2pf+qU2yWTSPtb/wDiHVTRNJLJJvOkK/zP+oUXm+XnBjdIcStFpX6MYyOvH0VGscBwDytl35yobFZLwnfiTfOATWuvOIGd8rYP5ijcFJX6rNYrnHGSKHOpzK6P6ldH9VBZLNVnboV0X1XQhNETAyR7qAqZ8gD2NbSh4r4dq+HYowxoZEyl5nFfDs9F8Oz0ULomNj18ab1atKxsm8VGS+Gj/Kvh4/ypji1ugkNLlMMl8PH+VfDx/lUNoYwMaDdcGhTQSMZIWm8C5u5fDx/lXw8f5UY5GB0E+zeGS6CP8q6CP8qFpjbSN2q8BGzSRsdIzEEtzC6GP8qLTCyh+VezzND7NNix7hkuiZ+VdEz8qNphbzLtto6vehBKxmmAwN3aC6NnonRuibdPchZrSA+yu6OUjLuKqGtp4LYHovabKDoxiWjNvgmwzhrZdzqYOWyPRGOSMU4jchFaxprJk2emz4oOaGuad4RY5jXNOYovabEXFrcbo2moRWmjH5X9x5LsrMsnDMKk49rsn3oGs3xQkicHt7kWSMD2HcVp/s15/wCWVorU3QTDOqwxCvOFyUZSMwcF+0N9ss33rBrDxCvwvDx+iuTRiRvejL9mymn3TlobbGbNL3jBBzSHDiFfoYpt0seBXPM9sg+8j2h4hc08H5d4V2aMPHetJ9nTmn3TyhFb4HQv40VYnh6v3bkn3keBWBba4+/B6uOrDJ2JMFSaJsnir32fanR/8OTFqu/aFlcwfex4tVYpWv7lfaNFJ248CsC21M79VyuyVgf2ZBRc7Ex/er32fa3RfI/EKltsZc37yLFakoB7LsFeDbr+2zArUkEw4SZ+q56N0XfmFrxxy96rYbXJD8jtZq/abJ7Qztwq7f0b+zJgttnqpHEVN44uV10oLuy3Er9msuib95Ph9FW22p83yM1Wrm42RBc00ynuyWs8RDg3NXqXndp2K52UA8Bmv2KylrfvZsAr1vtT5v8AhswaqRRtjHcrsQM7+DFrvFnbwZiVeDbz+07EqssrWq79n2YuH3r8Ar/2haXS/wDDZg1XYY2xjuVwc5J2GYla7vZmcG4uWq3W7RxKvSPDQjF9nwmR3bWk+0JjK77tpwVyJgY3gFru1jkwYkr/APxQfxn+iq0a5zkdiSi57g1vErQ2NhmlPctN9oyn/lNKDImCNvAIvleGN71zANks33rto+AWoKvOcjsSUcRgiyz86/K9uC9otz3NYer1j/RCOJgYwbgi5xoBvKMP2eLseTrS7LyRI15TtSuzKu3hXhVXG85P2eHitPO+7Dx/kEI4WhjByex2AaSfrP3MRe46W0O2pCtaRrfErSuN6uy0dZa77g3nc0dybFCKNH15BHFr2mTBrUZ5zftUmLnHctZ7W+JUj9K0tjxdRXuODB2Qmxxva52bnA5nkfM/du4qS32jppsu4Kr3taO8poEoN7AUTy3GOHUZ3lNa6RoldrOqVgQUScgrTbXdd2CxcAulb5KAMNWMaXJ5kfdc91cVqysPms1MfmA+iqSAsZWeqYG4kO4KS8dpvBdK0eOCwe0+BUcoOLCHehVbwosZW+qlia17zTAhhVnlJoOjeq1cBxLSsJWeqvtcNJHrNxUchIDusO9a0rB5p8Ljfa4U1RVNdQtfGatrheagW3jhXBtaLpAPHBOj0jK5tdXIp1ltDgJosKk5ha0rB5otvaQHcBVOns7ZBZwbwcRS4r05uzNoHAb1rB7fFhTopHsc07iV7HPIJbMejlrkq6ZlPxLpA78OK0thifrHWZdoELJ9oVaeq93804xse8NNKtFUWyA3TmHtKMtjlbNZTtQXsW+CD2zNFdzjQrpWu/DijJZo5GT8QzB3ih7REX2beK1uqNkbtIXitGrWZI3xYUZ7DaG2abew4Nciy0EQTNzqcCunYfAqjopHP3PYw1CIYNJBuEie6YGKVmcTt/gtIyJ7m/LQrTRGSxT9trCPVCG23XDdNFl5rVtDD5q5JC6cdzCq2B0gh7M1EPa4rnzsxCfFGL9DQG8MVffZ5oZd0kYx+i13e1Rd4uvCHPXSeq4Yq69unbwuErSfZ2nid2HDBftEIkA4HFRi6S85sdqkLGATN7nAqtmfKwfdzMJaiLU02dzczSoWq/SA8Gkq/DZ54Ze3E26rrrs0e7S4FOfNE9hA3CoVx8Uf4XP/AKq9A2eD8Ou30V20QOc3tsYf0RY1zi4ZtuFV9ikv9tguFfs8xEPZmNUNM1rj/wANaIwER9p4IV6Jrb/GKShWDHyt4Obj6hN08csBPaYtaxum77lF8FJ+f+6lvOk2jk6iJs8hYeJaCqNmZM7s6PFPviCz9k5lX7TaYie05v8AdaKCeW1SdmFoomzSS6CIf5bjeqqPcXA8MFpGhzX8aqptxaPnAQFlax7N8kjLo/VX57Wx7Oxcw/Vc9btHTqRNARbYGzXPvpX0TI7TadIR2f6qr4anjVUjtE0YHzf1Wjs1odaJOGjB+qparY2L5YmrWtWibvLQAtFZdNa5O95p9E60SSCzseNnMrnW6Z3aecVSF0kI4MeVeNue0fOAVhaNFZu26Ojj4Iv9oc6Q5vuiv1V60WmVx7N/E+iu2KDRRDru/qmutkhtMg3dUeSvNhDHcWYLVnmZ+/X9VoLDaZLRLv1Rdb4lMntdsMkw3XdUKslploO8NRhsrHWmXK85xITzaZTFDIamNuFUGaBhA4hat5n4XkK8bZMzgK1qibbaZWwHZjwr5oRiaW6N1afor02udzXOJJTXWVugps3BSivSc9M7ac5dE3yC1XSM8HlezWK0zEDpJCdVqNyebWzxzWtef+J5KdZbFGwHJ0jWpj53uMEeFTv7ggNCyg7lgy7+E0Re6edvBrZDiULVa3ye0HEa2LQtYOf+J5KdM6JjQ3uzT3VPOGgjH0V14DpXbZWMLPRYBzPwuIRs7Hyus0PSEvrig3XcB2nlYQs9FHZITdu6xuoEiscOse9yxaD4roW+QT3C+HHVaA8qIuDw67iL5ouib54okANA4KeX7x+GKiFMTitaNp8QuiA/DgrTDc5lhqNY5romnxxWq0DwCgIFdZWXhe/ksQCsYWeilkhiAfSme5RPETdZoOOK1WgeA5LVBTPFqEZ2ojdWswHxC1oGeinsssTSH68ZKq2Jv7o5NIwc7FiO8Jso6F+Dgg7BzTktaFh/dTbXZoW1ixdHTBwTJYmMAPAchaRUHcqtxhcdQ8O5CyWg6wwY4/osWg+Kc10DMd4GK9mtUbTC883Pd/VYcl14o7qv4KrdX9HBVGrINpi1o2u8QvarExjZRnGRqu/oiy7oZm7URzHJQ4hGayc3J2V7NbwSBheOYQewh7CrkkTfFuBCpO3TWbdOxuI8Qg9jg5p3jkuTMDu9aaxSF0fAIRWsaGXjuVaNeD5oyWBwhJzidsH+i0VqjNmm+bZPgeW/H+zzdpipM32qzdoYqgfcf2HoF7LrxlIzBwX/APugG8YSD+qox1H72OwI5KTRNf4rSfZ85Yew5CO3wFze0rl5pvZxyKtlebP8oxb6Ln4bzfvIsQqscHDkxj0b+3Hgq2O0e0Rdhy0dvs7rO/jRaSO4X9uPBy5mQWhnZkwd6q5O11nfwf8A1WGKo9ocOBCvwl1lfxYcFqPFtiG7etFb7OYXbw8YK9YbRojwYaj0XxLPyKTRxdc6zlWaS93ZBXQ4F3ZjX7LZtAztyq9brS+0ns1o1XYYmxjuHJdbWV/ZZit1kj78XLSyc48f5kpVyL9okyuxrdYYPqr8tbTL2pFQCgVSaDvVLNGZvmyaFW1zX/8AhswasSyFgWisERlfuctJ9oTljOwuZiAPaOfJV7g0d6/Zo7rPvZMlfkd7RN2n7lemkDEYPs2E/jWmt8hnk7O5BrGhrRuHJd2pDkxuJKra3aCH7lhxPiVo4WtY0bgqOdfl7DVcZWOH6KtL8vbPLoLIzTTb+y3xWntDtPae0cm+CpUVRih5yf6BGWdxu73FBkTad/HkJJoAjFZiYrIMHzdrwQiibdaEReFRjSqNlsh1cnPG9aSTCEHH5kGsF1oyA5HSSOutCFutIpGOhiP68jhpG1AqRVXGdAzL+q9qfnkxvDv5aMxnk1WBNYcZDrPPE8kh0jSWtrQFSWh2s4n6plHAyP1n48tlsnVZzj+SpIA71OGSAvLaCigZ5prWSNNBSnLan8Xnkq4gDvTGMdeN7crPKcmvG5asgrw38kjeIQZ2HFvJV7g3xUVpi1hk4gYJ4eaRSBUEgrwOHJFbouks5r5JkrcnCvJrva3xUr4Wk2ZxqHUyKfZrQ6gYKtP8kNe7XtYLiFpG/AzHWHYKqMRyOjtDm3HbinvhDnxsykpmE5lqdSSMVr2kDeuVyviiMclHsKFktZvQnopv5HlMdoe0cOIRnswfdZ1wKJxnNyWMVI4pr6loPaFEJI36O0N2ZWL2a2t0U3Vd1X8t2V7RLuLc06Szhzoh1TvT3u1JWDGMq9dc1p7QwRm+zpWsdvi6jv6LQzNME/Yd/LlOuGT8WYomIGSIdV29PM1YJWDFjlz0Z0fzCoV77OtDbRF9w936FaN4MM33b+THJF0T9FaP+CK/RUcNLGN0mCeZgYJGjYk3qssDmSfeMzHouYnZb4uyTSQK5jFL93JgeQiUNcz5kXWOYsl7MesEL1Hs7MhT3WhjoHtGTsj5qpjdDL241zcrLS3snVerlbknYfgeQidrHN+ZX/s6eRso6sesE0T3Hj5zin+1Q3aDJwqFsPsz+MTqj0WD2TD8rvQq7W67suwPJS0Bhb86Lvs6WZsm4RirV0j/AMytTH06Z5aS68aVVJJZPI0RdFo5v+a3H1XO2Z7e+PWCo+a4fmFEYrPzr/BXrS791zro9BitFYGmn/AZT6otm1L2NZHX3Ln5JHnjeRNnLHV+9bX6rnbMT3xGq51zovxsIWisbdK/tUNFpbSL3faHXWj90LRWaRzjwhbdCdeGiY/EulJc5VtBdM/tOKPssl2u57arnIBIOMbv6rnhJD+JhVyxtdJ890kLSSRhzxjftLsv3QnRtndO/hHqNUjo2CBkmcj6k+SLp62mQ5vkR9mldD3ZhYsjnHy6pVZ4JohxLcEGWRkgj3yBlT5ImGBrHHOWd2sUWe0OtE3Zj1WqV8PNNkFDITkiZBp5Dm+RcxI+DuacFnHOO/VKvWizyxjiMQhHZo5m2brPa3ErRwwMssY6zzUlFsk77RN2Gm6FJ7M0MMgobu4K9IBPMc3OC5ouh/AVqyMlHB4oi+ezPDRmWmoTQ2Cb2HfTC/5oMY2KzRjIbRV+1TvlduZWlfRO0IuaTUDIxuV+UB87s+5VaNEeMZoubnvjhKEXyWYFgzcx6ZKbM91kZkzIE96zjgb3axTpLTI+RrRU33YJ7ohooqXQxo3L2iVuu7ZBVbl13FuC5u0E90gqnPdAyRrcSWvovbfZy9jMGCuAWtIyEfIKlVkLpj85RZFQRR6oDVpHDUh/9yqYxXiMCuatDx3O1gi4xxytbiaOop7a2EPMnF2yteYRjhGP5qrgZTxkNVZ7OKADEhN4MWuxp8lzUz4+6tQiWaKanHVXMxscXazi52S5ye53RhVc3SO4vNU3IAOWYwPchfYHeIXNSPi8DgubfFL+IUU0ETY6nXN45LnLQR3RiircvO4uxU0e+mCY7rNNFE97Q80oa8VzTnxfhKcxkscrSKUkanfZ7XRsuV2lztoc7uZqqrWCvE5p0bxVrhRPY714heyTazmbN7eFqViPyGifG2dr2uFLsrE37OfIxlMnOFVztoe7ubqhVawV47+QzxDmXZ9yFmtGtAcq9VXmC5XfGaJ0XtF5p3SNqmWK0Stjb1ZS2tVzs8kndWgWoxo5HTWYa3Wj4q4aui3sctLEADvuYEIx6ckbr4rRRw2mX9myE4bVBz5nzg/Nh9FqMa3wHIXDm5e0N/iqVLf/AGlBsoENo4twV1tocKZXsaJrLTK72XLTMZVCTTOtLe92HoqMaG+A5KSsqe0M1pbM5z4/l/ohHbIgHfeAIGK0OI6pBvUTQ6WSWy9qMYquldO4ZtkOXkqNaGju5LkrA9vejLYJDG7skrQ26AOd2pGqjXuik3Y19E0aWWezbizNaznOlHVnOKo0ADu5C17Q4cCi+zk2eT5clSaP2qAb6VQjc59mk8UHxWp9psvyvQFoY9kv/Hx+q1aU7uUnR6N/aZgq2WX2mPsOWht1nksz+LcEJLLb3TQdkuoQm+12Z7HfeP1x6qsbg4d3JL+I8lHPq7sjEolkYszO3L/RaS1zvtTh1cqq5YYBZbP2qUWktkptD+G5XY2NYODRy3pZA1EWGz0Z99LgFp/tG2mQD6+CFm+zLPTcCAtJbpiwdnMrUj1u07PlvOIaO9aGwRG0yceqFW3Wi9cxcG7Le5CCzgPLRg1uSc8AxxuO0ckHSc/Lxdl7mis7PaJuDch4lCa2yl0QODG4NQDiG3cmBaCytc1h3NQktjtI77uuCoBQcOW4OdnOUbc0LRb30gGzC3JYXY42j0TobH5yLSSEsi3vO9COJt1v68pkldQIT2oGKxjYi7SDGANaMgFjrSnZYqmskjjgFffR1oOZ4cpJNAFoYqtsUZ1ndpNjjbdY3ADk9nhPMtzPaK00g5pv19yP7OgzO2UyFmTRyOIPOP1Wquajj6207x5TG3bmNwKNm84nlmObWmnop5eGHLMeDSnU7I5T+IKQ0yUTuLRytIwDyW+5aoaYHWapbM7frN5YvtCLNp1kyVmy4V5b7Rzkf1CbIw0c01TJmnPMcDyaSPC0R4tKuSYTx4OHKWuF5pzCq3GF2yULNaHc31XcEMc0YpRXgd4QsdtNWf5U3H3DJFqT/Rywqxzc2lUrcm3sTopAHgjFpXMgz2J2Nze1X4nVH6cpjlaHtKM1mJfGPUJsVq12cd4VQRLG5GSwy6InIdV3ceBWgtTPZrRwdkfD3C4DRS9pqBBJj4jEFaK0gRP31yK0lbgzZaYzi3xX7QPabPuni/mr0Tw8ctyVge3gVpLBKWHsEp1m+0IS5tKVIV2Xp25SjBxVTILXZvm2gqXtG/sv9yuj0T+0xF0EntEPZ3rQWmKjD1HDJX7FaLnyHFqbHa23C7J7clejcHju5bssbZB8wRdZJXWd3DMK5NFpYBvbrBAx3rJLnzf9F8efRWhrOdkEhFPNH2q0ezg5QtzK/ZLP/wCpIrtrlMMR612oQlYRaHdtxr7hMj/IJzYBom7nrTT1tFrG0NpObGwWaIjC9mq/aD5Azi0Vav2YMu8W8tXENHEq5ANK/cdyraXYdhxoEI7FFWSlLrG71R8ogGdzj4qttieX9twqxAxua5vy8tHG9IcmNzK595gZ9xFjIfHgmxMbFZbO11XtJq53ohB9lREkjapktJNPpJjmChG+A2U73nEHzVWkEcRyFzjdaN5RjsOrENq0OyCfog+0v683HzQa+6IW6uiiFfqtFDVsXAbkx9RM4ZtdgCgyaM2bx2fVVaaju5KuxedlnFe3farxHGMWxE0C/ZYaxt/zH6rAp2mkx6t0UaCi5zie087k6Szhstd0mfkVdlBs7+D/AOqw5PYbIeaHSSJsLT5DFxTpLos0Q60mfopIGlxLndIeCq+ohbtFBkQbNEOrk5XHVif2X4cjpDtZNHenWyfppcceCuxAzP4MUk0sggaBgyPFx81GZMLjbtEXOJa2PGo7SxAtDeIwcrtbr+y7A8kUObIR9VrENA4qlnjMvzHBq07pucDhdYzAKWU5lOe2R0J7t652PSt7cX9FqPx4b1aPwFSeQWu7HhvXNR6Fnakz9FEb75XPdR14/wAlKKJsjZ3MkBu0OIXPRVHbjx+iqx4cmS9ktegVcZWWTssxWs4WdnBuLlBOyprquLjVaWI6wyUcsUxa/JzXawqv2iItHbZiE9gIeHDcprDJmw1aqucAO9Us8Zl+bJq5+XDsR4BNlibSM7uCfGw82/aFUyazTVB/y5MfqqTxmH5s2+qb9p2PEf5gamSsOBVXvDVzEV0duTD6KtpeZ+47Por8fQu+igZLrxR5Y4pstmlEzD1JM/Vez2xuhc7Zv8e4oWS2G9Eeim5Ltb7+wzErACzM78XJ2lBlc7Nz80JYidHXB43ISTipyvx4OCoS21N4HBy0tjebPaew/C+jDK3Q2lubHKpKuwtM7vky9VryaBvZjz9UWGPPrb0ZLM8ui48EdNeaHZuYqStbbYtzm4PaqMebXZh1XdIzyV6J9e7eFWR4aO9Us0JI7cmAX7TKZB2G4NV0xhtMnNzCdHFKZrOc9+CxvRD5MvRaaDUk7UG/xatHav8AqMy81eY4ObxC1n63ZGJXNRiBvakz9EHzuNof8/8ARVu6N/bZgsH+0Qt3UxXOtMbuIQuO08PqgCdE/g5ZiiuR1nk7MeK1nCys4Mxcr128/tuxKq2sZ+TBF4eLU3cCMQqOvwPHBc63TN7Ua1JBXgVrPa3xKpZYzOe1k31X7RNRv3cWAVI2BoWStslom0bDO8tDcTSqDo4tftuxPLfiJgf2ozRa7W2pnEarkW3JNIOrRbYsreGbiuZic4u67sVetb7vgalczEAe1v5b8dYZO1Hgi51y0MG/ZKLYLM9024ZhaX7StWib9wxaOxQaFp61KuKElpJY08dpUijAPa3nlvxEwP4x4K9No52ca3XIMsMBZXae7cjJa7TekOYacfVGKzNFni+XehJNWJnftFBkTLo48eSlFegc6zu+TL0TRNo5q9k0KDnsuWXcCaD+6raZL4GTMm+i0cR0UI3BXujh3v4rRxNoOShFVege6B3y5ei0LtFM89nCiNqtV0SuyLsS3yWntb77G41kNSUYYebgH1VxmDBtO4IRxijf15KEAjvVbPK6H5c2+id9nxljnk0vxpkWkETTi8x5nzRutDeLkYIjzI+qbEzM/RNhZkPryUe0OHeibPMYx2XYtQbqFsP5UPaJTJTqN1Wq61oaOAQszDqx5+KwxUcfWzd48lHtDvFPkhtBa1ordk1gn2lkjWPe6r3EVV6Qmd/F/wDTks8P7xQ+Y/8A9uUffjyazceO9OItTjDgCx4qnuZaCyCuy0Y+qq1ut2jieSE/OpKnAqZvB/JeLaP7TcCucmdLG4EC8MQopJp3yNI2MgrrGho7uSZu8C8Ex2/JSWYnbxHJeFY39qM0KjtIlc59duiZK5xtFRUF/K+J3WTo34EIRPPMv+i4hP0JMLz2cj5L2d0z2WZ52mq+Bed23Ynlcx4q12YVM4zsuQoaxb2oGJzScxXcVcDnR03A4L2O2SyCMaoxoFzbQB3cpa4XmncjNAL0W9vZQezLe1Y0J3tK09ne5srMm1Wi+0DIXHZLzghdAA7vcMlmox/Y3FUo5hGbCrkzRf780bRZJH3XZ0OSuWpt20duTFYe4XNGil4gZq8Wubwe3IrR26MVy0gTBY5XyxPyFVopI/Z5vm3+aw9zXZdd225oyQVkbxZn6K7aI9bttGKD8Zo+yShHd9nf2SsMfcIljDq796v2J9D2XFaO0wODtzhgVebdtPySZq68aB/Byq01HdyzfjPLU4BERc+8dlUlm0UZ6jEYrPHV+4sNVftclK9Vuauwxhg9ypWjh5+XgEXTvuxjqDIKtlqX3aXgUJJSWMPWchdZek7bs/d0Vnbp5u7IL2n7Slw3Rr2eFo0tcSFveeO4IPk56XvyHu+z2JumnOFRkEx9rfpbTK7LsjehHHQuGAaFeeSa5NQltYoN0f8AVAAUA3D3PZrJzloOGG5RG0c7OayO7lfkN0K63ViG5XW4MG0/ghHG2jR7ns1nxnfw3KWR+tKNXw5DZIHfjKoBUlVd0z9r3BZ4zzkmfcEztv1nHkfLvyb4oudiSg4jUi1j47vcbA3amdTyUbeWQbmaqgjoOJ//AKijbwHLG3tSNX7x5YhmdInCn0/srWwmmIOPLXsmqkj+7eRy0KtNnGVdVRyjNrk0gjWF4ckjN+YT7K/ajOHh7gtAwcMDyezyHnG5d6N1wNMDRV6zTgUbDaMHtwbX9PcdFIMD9E6J2NN6FcYyhLfAaeKc3DnGXmvHFexW3AdV/uunswxzMaD2G64K5JqyBOinpdk1o3cChFaKzWTdJwQfG6808PcpI3W3PGYVc29WRqdZrSdVwpf4JrtXS02mrQynTQ/or0Tq928e4WuAcDuKL7MbjuwckWtbeDDVzc6K5aGhsm471WF/tVn7J3K6Dck7J90346P7bc0ZITpYxvGa52PDe8qtml0kY6j0RO0wPGYKDmODmnePcuvaHt4FEwHRHs0wTWzNFzi81Hqi6GR7R2XbKaLSy4Tvbitoqb8ZVZHjw3qTVDYqapKa99+X5Yxgqi41pGy4EFGO2ukgHVZeN0+aAiaA3u9zFEN5x/dkmxyzBgJ2Wp0VlidJJXhUK/JI2/8AdjJNbMwstX/FyPh7vOPF7s71n7PDw4o3Wh07Rid1e5FsQOj39ya4ETEbTcqoQMZ7M8f5TsD7hklddaFdjd7PZe1vcm6O7CK4l2L3Jz4dt+GPVCvnY60hWlZELSP4gtR2sM2nAj3PY7BrPOBeEcPabYdqnV806Z79I6l3RMGARxpHuC0ktWw/qrmiEkHbjGPmFejeHDu5brNad2yE63Ww85ta25FsAo4gyPmeMB4cVLFGXy3v8125EmpJQtEhLJTizuVLUzV+9Zl5q80hwO8cj5X5NCdaJcnHBC8cdzBmVJNMTZYdzG7TlEwgtZHlXeqphjkMc7sXcCgy0t0Tu11Ty0zZDq+apwWjs7dNJvpkPEpk75b9ovarRg0K87acalSOjFXNwH/9VNNnkx3sfkVo5WmGXsu3+HJZW/PX6Jnmi57g1vEqkA0MX3rxifAKzXSTerfLzmjll3f1TI8NE94DhxXNHTR/dvOI8CqDVeM2OzCkbxCtEfbaH8l3bkOTG4lc87Qx/dsOJ8So3sAbE4ZI5fRCGd1RdpGQcWrXHtEXabtDyV5jg4Jlpb0bjj4IEZFVJortkbf/AOIdkK/OdPJxdkPBOHVOIV+J1143ojSaK0jG+Ot4p1ntguFwwlbs/wBk23WfpW7V1Y9M3aHJekcAtX9mh4naP9E6IsqHZk5osds9V3FBjX6oNaK9G7Q2hvUOyVobS32efqP3eq9jtuz1XqvJcbWWbsMVbS64z7pn8ytHdDKbJbuVDVpGTgqvOlb2CEY+mbvhlz8inS2Ml0X+ZA/aCqw0dvacxyVJoFcsbNId8h2QtJaHaaTvyHkqjm5e0EWVLQfGipOzTjtUxWkskhZJ2CtHahceOtuVQaju5KvdjuaMytatng7I2irrGgBXhzcvaCDC91wHbbjVXnR4cW4KldMzsnaWo6juyc+XRtrLL2Gqtodcj+6Z/NXAwXeCLojcfwJNFV1csA1uqgHAsB3IX9U8VVrgR3clSUY7IzTO7XVCv2p+mdw6oV0tBbwTdDzfdmF0/wBFaomG7dkcNXxRua1M8U2SQm9vbIAVzUTWeA5C17Q5vAqtkfej+5ky8itHJWCbsSKu5YG+foi1pqOAyTS46SvUa7FVn1R2MCfVXYo2xjuHIWvaHt71zDtNF9084jwKoXaOQZsfgVfe8Nartkbqb5DhRYE2mXtuyC13aRx4FB1pqxu5gKusaGN7uSj214HeFvtcH8Y/qtWQV7LsCqDXk4cF7RaHXIh1jl5BaOyg8DMVjrO44oS2mrY9za4lBrRRo3cl7YkGT24EKlobpovvWDHzCLmzMoO9ezWaojOGWLlrHQM61Dru89yNmso0cYzICy+hQmnFIeGOsgAKDk0kbjDL2mKlrZq/esyRkY8SOOy0FG1SM9onOy3cPFaS1P0pGTeoE6GHhRx/ksvotLIOZZ3bR5S+yu0LuHVPkrtrYYj2hi0plmjeNCMXO3Ix2Ruii2RM4bu4J9oc4yOcdp2aFnadRua/+k2o1I9Z3IQRUKtlfQfdO2f7J2maYZQNl2/zTpZaumk1gxoqSg+c6KJ2Iib/ADKusaGtG4KOHsiqLzTD8KblrP7v6cl17Q4Lmjp4vu3nEeBUDQHMcypc1wpRRx2aMvcBi92DQhJO7Ty9+Q8ByWU1pnvQ1sxne/sonA9Yb/7cmsNYZOGYWuPaYh1m7QUNqFdGatyxWqDZouJ2j/RagxObjmeQuGbMUDjq4b1HIOqe9MkaahwqnSwnRT0wc3f4oNtEOt1ZY8v7IWbROlmZgKcFetTrw+6bs/3VAKDkN0c4zELf9U2VubfFNtDaatKhF1ldo65xnZK07IjFxZmCv2aK4PvJN3ktI8mWXtu5TG/913Ap0UgoR4oPZUOCuSAV3tci1nOMGTHZjwKMFoa5zBlhiFn7PCdzdoqjG05THK2oWIvRnJwCD2Va4b6IR2gXZRk7f5L2iB1R22D9UyPQVnPfgr1rfUfdN2UABQd3KWStD2ncUXwc5HwpiFvaVctQrwkGYVWnTWc5UyRjs7GxcXONaLSOJklOb35+4WuFQdxRfZqRnsEYLFro5O+gC5zaHXbmFWntTabWRXSCGLgzaWq2nf7lHCoR0QbET8oRc0OuDrEraKFyJrncaoOtMtWfdsyQDQGju922T2l9b073BjfxLUY1vgPeLXN0zv0T+ec9vZrgFcFX44BqbJaKwu7jiqRtp37/AHanJaGFmnl7Q3IPtLnkjqAq7sR9huS5qPRR73lxWpVz97nGvulziA0b1ds7MRnIjabSw4ZNO9UIpEOohHFFUncKoSTUfN9B7rnyEBoT5IYbsQTZqC+4VLijFDscVs/RCa0NpFuaRtIAYD3HPf6cU1z2ARvfuQYxoa0bgtFEedd9FimxtGG80GATYoxRo9wjAvfgAnPlZWgBFeQNeRpaUCLnGpKrwQLhzkmsfcgs7dp7qpoNLxG0AgByTvrhewxTuc1T1aptZLzWtrdBy9xoYaUjqoB8g5bLR1w1OKaTKSdxqcEwl971TDxHLpGvNxrw+6geWSPtCikhJxHiv7FOs5zjxHIWAUbwTX1Jjcbp93SsGo/9V/ZCOTonEeqruKk4jFGGbonH/wDj7u4St2XIse0tcMxRCSM4oEbW8KMMweWkr2a01uZAncqj6e4WSNDmHcUZI6vh8MlhgVoLRiDheKdMzMO3IQWvA5CQqoPp7pfHSKXwwKuSsLStatw7hRaeyP0Uldiq0VrGjkyvFYGvh7tyVgeO9F9mN8dg5otdfZKO8Jr66CXtsOB8VS0gU+9bkqtdeHd7tHCoV6LmX92S2Hf8yuCpex7igH58Qqtde9yb8Z/XlzpyZ33dkLA0b2WptXsunqNer2vZYj89SVzbNbe85+7UnBa7qv7AVXHQWbgN6GiLO+tbxQihBo7qBzqIPtOu/sA4KgFB7tXnW3NGZRA1IR1VdAvz94wV5/pQrUF1m95V2MY73HM+6ZJDT+aDHO0cVcGlPibQVGaEMd4QtFMs1kfRC0Tise5vFcPcdJIaNC3iIZDgFZLPEQHsfWiO95yCL34uKoB9E26Q5zsS4e4XOwA4oyGugZkp2jK61M0jw0u2Wnei1p5tmC/+lE2XCIGrzwVRl7k0mbGajVF+HktVx2LGmh3HwWf8Sijv4V+8qE5j350AN68B5+5P8sQCjHcOQucaAKFrCRdJxdVtRxUZvg/+o4ppvA/+o4qFlaaoF7dXhy07TCrO/wCXlvSOuhX2EFr8cFh/NRuJow4FaMG6TsE5P8ESg+mttIA7ceqfcdZGN0sx3Dq95TmObRwzFF/ZaKZ9x7Os7BSRPaYidmvWCvNHONy717JLtt2fd/ZW3pW7Um7wRa5pDhmKISR17xTNQWj5S2h4qjmiK09X5l7Laa3NzjuVR7hvbO+qe6wjmxvOVe5FrmEOG4tQZJV0Xhkg9hAkIqGjehFLWSH9PBB8bg5vuu9pDbg3ncnyQV0fVvjFy2S1w3FoQa9rnSdrAURh02kHZOQWrqu3g+8TaAA7cRtIvZq8GOpUosuvZJvbIRRc2/RupsVq0ptIxfa6j8ULjtbs+7Q4hVYTHM7JkY2k54wl3Nqhfq1x71zw81G+MaSzHaIXWU34zyHG87gFcL9FBXEhFoDmWZraB5OPmhcZpW77jgr5e9lc2VC9osoFd8bsii3o5RtRuzHum87W7Kp/lg5BSyyFlerpZFdsrXB/yyoS2lzpJOzeqF7RZDopd46rvFaKQaG0DNh/l7r2QEOcM3nIIuqZHnfvKcwlgveVEGM13n5ihJML83jgEZ7IbknWZ1XoxuGinGcbvcq7F5yYtPaHgRbv6BUs7L8gyO5qayV97jUHFBrRVx3UK0kgDp/0RlsmG90J2XIjYlG1G7Mcpe40aMyhFHUQjIEfVGOzUaOvP/RFtlacHdLmSU3SEvIFMWqgbj+BXntGmfnhl3K/ZdjfCcvJauDhmw5jlbYotp+1RNbvzKtXszNIR1zsiiYGuMk78XSnNEmtT3Ku4dwRleNab9Ffs2vFvhP8lVhyzBzHJLJvAw8VfdmcVE6VwY27XFc4DDZOxvd4rRM1Y2Cl1q3+RCYNbV+ZtVaHPBfpHUN8g/ouarNZ/u+s3wV+N14cltd3tCC1sXHJozK0lrwZ1YBl5qIg3eb3PuqLXJofvg5bdfG0Aq0RPAe2uRxWFZ7Nw6zP6oPjcHNPBQ8LpT4/u3kcmihbpZuG4eK0sztLMd+4eCnF5t6/XGTH0TXVxHF6/wDkjA/W0Zy7k+Ce9NCBXS72+KZvBCuHCKXDkqckWWbVj3zf0VGDxO8r2lo7nLd6oio+q9mtJ0kT8q7lSSstn7e9vim26ynDPBB3XGDhyF73BrRvKwrDZePWegxjbrRuCM8TRphmO0sh6FU/kUGTc5D+iD3G+3dNw8ULNaDzfVdwVRyXpHU/mr01YrPui3u8UGtFAq0DZhk5GORtHD5UMxTg1XZmmSI8UJoH1gPAfqhSrX9l3LTbkOyxuZQltePZiGTeTnGi/ufvWIvM7TWIMlFwdpkWKvtvmHc6lEBIa96Dm0LTv5dDANLPw4eK01odpZvo3w5KSxh3ei6GksfDRi8FzLZdLvqyio8XSNyAk1+/eqtdXlMNlGkk3u3NWkedJMc3nk1mh3inmtWnqUTpIw6HddcujU9XVdfOHmjjcYrrK0/VNNqhledwa2oC15Gui+70YVI2Bg7hyh3Rytye3MIQ23DszDIqqvOdQIiPV71o46uruTTdmNq7g0haS0vfG3gQKlXY2hvLjqvGy8ZhCG25ZNnGR8VUfRXpHABOD6wx1wY04uRAoGjdWgWoHA7zpAhdviPe+9krrMTvcc+XHVeNl7cwhDbf3Ztx8VUGoRYwtdPwJyRtVrLscm3sX/2VSWtaMm1oAsKD/wBRBjNZxyAer78ZznjWnKHgmOVuzI3MIQ2wXTulGy5Xq4LQROGgGZ4q8+scJ9Xr2WAtYxuB/oup6lZt9ShapAKdTl0jDophk9q0NrGjk3O6rk6Ynw71Jb7URSuHeVr1gs/Z6zk7ANjATpDTHLDILd6KKEUocXEDcgBgByaWJ2imHWG/xWhtI0U30d4Kz2RvWN4oQM5ydwwaEZLQ7SSBtANzfBCm5tVK/wCbsqtMP+TeUj6VHdDfCZ82OVOTTWd2im38HeK0U40M3ZO/wVrdjjKmwWfnJTRteq3xWlkOlnObz/LkioHHU6rA5RktkGPWiDUdWb/otCnZjlv5K2SjDdvPbucjUaOVrMWO8VaWPN1pAfirtn1Id83HwV1g8Tx5Ktv0e3JlP5qSE3weAout9FHWt12qaq0upq1uoyWXziORWkZVk7NphzTZZXUcNUjfVXpqxwbot58UABQchY4VacE6PHux3Lf+Zb/zLRydI3PvTnwC9GdqHj4LSwkuiObSU0tfpHOya3NCW1ZdWHcPcNphB+doK/8Amv8A5q4+hgO6taLT2fXhPVG5CGcjRbiTsrR2fn5TkG5LT2k6SXdwb4e5deKHc4K7IMNzr+a6v51eY5pac2VqtPZq3x/l3sWoMtD2Mk4g5rRWMX373nJqL3HSSnN59wtcKg7lfso8WEoskaxw3sc4oSxSNx3NOSAcbv6FX5HXDw4q5Zuai3yf0VGjHeePu3nNpJ2giJYonM+9FahakgkbxahR1CtcVPciyOsMG928oNY2g9269oc3vXRBWwuP+c/9UGMBNcmhH2pjXO3Oa4q4wUHr7xDwC3vVIbQTDuYcUXvJQDnXRX0WjgbC+mcpaU1xY18w63vFrheaUILHNfHZOIYqvcJ5u1TBvgqyvIrvzQaCzD/gps090RdnR0JQZG0MaNw90hwvDgUYbLaHXPWncr9oOmlOLWEfqi6dx8gtp3/TCDI77nH5Aqu15j1qZe65rwC3vUlns80mgyQnlN6MZDitBEdfu3LN/wBF/mfRY3xE3aOCAAoB7jhIAW96MYkfoA7VqUJX65zbXq8nszK8XUK635l1/wAydaHbcuXh7hEratTnkvLdhrisMTvccymtORTyB8oCy/iThcOIzEhRbcJJOYlLVG3gOUXsm4qOItdzkm0mRtbdaDXlgN0O1d5og0RNb3h5KpoYh++UGi7RwOXIZN7hRON3WbiCgXi7dAwO9UAoOVz7jXmPWo5A3GNHZGSOrGPALqqOXec/HkM5aLzMapglYLr9n3b7RWSPHxC6v5V1fypsrKVHcmyNyKE4GLsCrsoFHYB3D3jaIQNEcwG5L/4L/wCKuSGsR+ivRCge2taIslGo47fBdywWvi7u5SyRt4LMviOTg1b/AMqvtJa5Xmx6GTjd1Xr2e0sutrnwQc0gtO8e993J2wi114tPWGR5OeiOgO4oU5yLh1mqrSCPfdonmInd1SgJGEY4HcUHSNLQVeBVH4d6q01961OklLI3TO1bveqQxgd+/wB7gqVvFVrdaqxRue3e6iuwxzF53UCbJa/+mEGsaGtG4e8XvcA0cU8R1ggHX6zvBfs8fNDaxzXNxPad9XBBjI3PcdwTZZ9ebsnIe8STdXs1jxrgXjer+pJaBnefQNVWsDePOXl/dCONl5x+ZcZTtO942Wzur23D9FdyaNpyfDUXi7UCLnuDnHM1XU9U2KMMLj3psUYoN/f7osrDrv2u4ItywqUztN1SE55z3Jz3FpccV1PRRQtu6xxIG5NY0Ua0UHuPoaOfqhYbW2mvGThVNUUNe9Zj8iwLSf8AlUKgZVuLhgYP5+5KflKsjs6GuSby2el4ap2WXkKmQjvguramp3QBQHW2t7acjUQNp2qFZ65EmM+45p3iivHTOLDSrmiia7nT4ZLrqSzmutrCvJHAOsau8FebnHlTgo5OtkfH3bzL2jfldXXXWVx9dE/6FNadiMV81ebsOy7loJemZvO8e6WkVBV9gc6B2+9kt/qv7r2e0tDoTkTuV9mtAcu5Cz2jotzidlVrUcl6OPSHeKoHkLXi805hGWAF8O/HZWX1VHNvN4aQhc7cYBsu0lSrrhfgJ3nDyV+N4I94skbeaeKMllF9vYJxCo9jXdxcUHMdHGOzfRIN3vQvEMP0PJUGo90te0OadxV6zNa75HotNyAtzaSroIJHArArX1XLuV2utw5Zvxn9fdjjOuXHG7uTtfEbgrjMG9y5xwqcqlXLsc1cmtlUcM7fZr2WsaFUiZic3HP3i52e4KNx1ZX4CM71fnuvo7ZGy1aQTQvrmxzlg2zsHdVNlLIxATQyUNAgYWguIxfx968/VHFPhv3WV3fzVWTxtmIrfcFT9n8RGtqP8iEcV17zuDU5l27ax0gOfvGzwO505ngsdYn6J4h6oqcMSjI95qfkyW0f+mto/kTX2iOjZspabPj7r5X5Dgn2iSrsa0KMkpoTiVI6bmdKbwBVwXrjOA3rr+izf6KZ8EeklHa4K83PItOYPuRWcVux4nkmikN1jddteCdaH0jszcKOzPetMy9dQwlPgo4yJq9l5xUAc20XjstldghBa6CU7Lxk/l0bdp/DgrO0g0u44/qhE7aiN3k9msrqXcXy7h3KJkd57420JY67iqmOYD5pqhV0UpFM9PRCS4RdNduqbamtrZ8nx9Yd6ZLG4ObxC+WIfVcG3gUxx2snDv5fZrNjOczuYOKmgcNM7O++W79E6MtvEfPRZD8yjlFKtPaT4Wv0Tq0B4hFlodec4XY3neq7sin2V1A1+WO/3BFEL9ofst/mnvN6cuxfXceKqA2h711fVdT1UbLodIML3ctBaDVsnRy8UHto17TUFNkaces3gfddZovhx0kv8gqGhjOy4rONf5afG+7K2mqEaACUZNKFntDxo9x7KqMRyhpa4g9bk9lsuMh23bmIGCmmGd7rIsfca4Zi6qjRHxars8sVynRtaU8NIhbndyqmtkdrcVh7tTrPODWDMp81raDI/qjJqMjSHR/hyV18jGDiI0GQOveS9nkvGzkbQzCuXhLC7Fp4qrTQ9k5+6XvN1oQmlbds42GdrxXMFsR/DVXZXOc7uYrwVYsV7ZA4h3XYc2/2Q0v5gukb6qb8Z5bznURazUHdmVeZzlqOXyf3T5ZJDedtVOC5u0Rsd8yBAs5j+8Maq2Nt/tURY8f2QstsNfu5u14+5gjTF3FOJee4cU2e11azcAEfZ7TUHcYVjLUn/hJstpdebuju0Vy6LvBVbWSxHNu+Pw7kHscHNORHuVetHGf7IyWvTR8KR1qrummuDIaKi25v+mmxxulqfkVK35N7yhLE7R2huy8IwzN0Vpbm3j4e5cYCZ3cNyze6Z+QcnQQ67/8ANeP0WzLXuX/iF/nrSyaTRM3O3osc2rThQq6+r7Gcnb4/7IEGo5RZ463GGmBzKEj+ij/icjarVqgbEXD+6MkrS7gKrYf+ZbD/AMyycCeJQcRR8msV7RZtWbeNz+4o4XJG4OYcxyOecgKq0WtwxccFeebrWjNCaRtIG7DT1lFGMQBUiq6P+JdAHf8Aq0QaIhQdQyfzUNbKxpvDW096iuPH9kLPajiejl7X9+S0nAtZSMB31UOA1Wcckx2TZG080+Cx4025B+gV6MUaG0T6xwux676InQ2Ud7ZcUKxWUnjJJQrZg/dcp8ASH4BvejI3nGuxki/otIDUvN4qvFqu9WVgkHjv5BZ7PrTu/hHErDWecXPObiopiyE11SZslTmXA7mZLOD91f5a2mDwV2TEjAnv4r2W07fVd2wmzNwcw7RUcwNbw5A1gvzPwYxGSQ3537Tv5JzHCrSKFPgdSmbCRuW1H+VbUf5VtM/KjZZSHxvyWhmNQcIpj+hRvGkRN1wog5hvNO/kqcAjFCSyyDakHW7ggxgutG4IxSCtfojHI4dxu5rpB+RdJ/ArzX63giW0baRmO0hZ55LzMgbuysMRy+y2Q6/Xk7Cutz3k5nkw1JdzqIxyucCPkV5srgfwKtotDxKMiIUC6teJFKhBrzgqsy5e3I7BrBmV7Tadac5Dc3w5dJA7RO4bijG58zO66i2k0zjxjVRUxnjuQFcQrsv5lUG8OQySOoAhNMLtnGxHx7ysuTEIvE8tOyKK5oZvxFi0kOD+5Y4LaVqDDrMlc0jzVSaIti1jxRfI5BrRUnIICdw0pzwqrlktN8nJuhwCv2qQTO4XaAKgFBylkgqCm2W1msZ6OY/oeS844ItjwRANe9aW1MlApq0jqrkVotOj/wCWgxjpy4/KqveZZOJ3cuKM1mF6A4vh/mEHxuvNKwWuiGlae0RT3c2GMLE2st7ysrShGwWjHedyutJc45udygg6OVuzIMwvZrULloHo/vHJg2/IdlqvODzI47yjDFzlpdtP7IXRSfmXRS/nXRSfnTYxG8De69kmxswa3koRUKoq+xnd93/ZBzTUHeEQ3GV+AWmfquOW9NnnFKbEfZ/utA0BzRicV0Q/OuiH510TafjTGXebbiVQZcgngOjtDd+53cUWuFyZu0w7loxS9KbqiD6NA13IPeLtmGyztKildRhFaDFbMfqidHZnfienG7AQN0rqKPmrM2mNYTU8kcFKRnWc5ez2s3h/ly8e4oXrt6R1TeQ2cGea0EGAadaUbkGtFArTIDqHq96fjZs+ujjYfLNYusg/5oxW1Zv3ArSzUOTsOQzQCrDtx8U2RjsKqAt2on08loINe0uyHDvKe5zy+R41id55H0pebrCoqmv00DjwjbRDnI2913FdIz8q6RvojEXikn6qhwOYcNxTrPPhO0fmHFSWOR+eLQqnWecGt3kozzG9O/8AhHDlvs6WLEKpku/urpv4V0v8Krpf4UYpNd2Tgf1WjeSWdST+q9kmkrXYw+ivON0cSrrassY3/ef2Qa0UA3DlLDqv6ruCdFI9wcPlXSv/ACrpH/lWkY52kHcr0R0doG23tLQyyPeyuZbsqoy4o2WynW68nZQa0eJ4+4WOwO5w3K698hG5wCqHy+iu2mWckbJu1VHAt7jghV2qqtzV1vOTHZYF7RaNec/w+6WvHmM1eY6V7O0xftHtTz6oyNjkbFuLhRUO0u5GR5u0QnnwgGxH7xaaiu8YIyM085/FVOlED43DiM1kVNaLPJo5dIb3A4qlcES4ru3BB3tdy0HsxVTXSWt7YeFwAlUY2nvOY8VBToZecibsvP6I40arjD5rSWgTtGbNGytVQzWsjvasJJ42DNzxRBjKn5jmfedaLJ4ujG9Oe9tCOtuKJJw3BX5WSPiGejCpS2XRkCVsWpNjYy0Di4nAK4ypO9zvdocHDZcMwjDaGaY9Wm9Pe+NwkpXawARLdeaTZH81V0T3POZvZr4d/wCdfDv/ADqgs7q/jWXOOxd7pls+MGZjO5OmfHgMgChNMNVmyNyc4bW4IudE0k77y6Fn5l0LPzLo2sPcUZ3No+T9PcEkJ0czMnKFkzADHmE6+LsEfV48kj+yFsxeq2YfVE6Oy+IOsi67ZHV++OKkddgFG/5HIxFrhVMs0rhJFXVLs1oIqNvNxfvog1ow5JY9+afr2YY9YIjSWH0xWMllb/zW4rpbMfwBSNvMN6M5crpbPhXaZxT4omVfKagnci95vyv2nFN5CDkVLC+0QMumlwsxTm6VrBxIqunYf3V0zfRBwmFRjkmStNQ4LSMwkZkVHaq3ZGnHvXtU5vPOXBoQ7vcvswikxC+I/gXxH8K6f+FNkEteIpmqbTTiCi28WAYhaOaa8xgxbleQAFB7uqbkrcnJzHyPa5uYurpn/lXSv/Kg+N5v8VehfoZ+u0dbvTYPan3K43m5IaPEHG9x94seKgq9pZHRHIgLpZfRa8kr3N2bwXcgATQ/RGVz9JIcid3v4p0sDnNd2AcEYbR7Td3tRuVpXBVK4jgg05KrTX38S5h4sNF0kn5la6/fO/VUqKpl11470x9nF26ek3BVlfp5e0R796uCux58VV5RzxGFORrNLLhgAE2a0SyBuYjO9UGA97ijxQIBO+4E6oI7ijQvp8q/8QhGzTDi45BCNlTxccz7znyYMG9X8WxjIL2iRpDLl267rFGR2ZWw8+a6J/quhf6r2qVpDuoD+vvCzM2nYu8FQNLiMTRMLMqK60Xo4/1XRfVdCPVdCKeKjhYNWqaxuTRQe49/6q0WomngnRPF2TPHkawUq92/gtlnqqBsfqqubGCcrrqoatnPe5ynqGgl9NXLkA5IYmnI4kJ16rmbJceWaQ9UJ2MIx6yJv2X8yBvQj/mLbs5/CosWY1GHhy6KPGV30UEoPrxVRtbxwQKB5L1+KMPbXnEW3mOHy5LpYvJdIxdI1Ps5eD1mrRtF+V2TQtHL1xgQvZ5TQtyXcfcfH1s2nvTo3O0bmZ1C6cei6cei6T6LRvdzbsu4qWe7Ro1U20RmhamysNa5jh72liN2Vv1RBmII+VdMfRZ1THOlMQHWArRVs0l+RoqcKVWgnJ0P/tQcw3mnf7xa4VadxTponu0XCmS2yfLkvRyvfL2SxOfkeCAlVRlx9+jxjucM1Ugvj7QXOGUH5QiKOucSKIUVQVQ6p/2FriY5rXaV1S45YqsdpgmlOQpeQkt7mEDKNjaINY0NaNw9/Xz4IgGjVePqjW0tgHhUrQtt1Y+FyiEcLtI88Ar8p0kv0Hv4q6w54Ivea1w8EXQ26VrzmGsRc6Z7jxIWDyFcjmkpvdTJCNmPed/vEvwA3rRRFwhGXevaJ8IG404rASNYMA2iyesdKsp1XnRGzE3lQZe6+V+TQpJ31vOK1hruxKl0dTpTRrRuWw5dE9dBJ6qujcx/eU+1OFDstr7mJojToq0HzKzRUz5xyBabkg2XLRS6kzd3FCO5eEbV0H1Xwek/eTYxZtE7sVQ//FsP/qKPVuVqbvDkcjDF+8/goGhowBNVPeFQ5yDJMYDk7s8kxORyTqWeJ+PWKP7BZ/G8sLPFIfnOSxs0DfwuUB0bBrhHxWji1pT9ESdZ5zcphTZNQo5oyGyU9VQi48ZtRbw5I5Qxj3NdTXyTXlkLP+WUCGQ04nNZRLKNRyi7qlaRmN/Wqr42mGoUctBo5NqqBFZouG8IPaa+4LZGNV2D1evRAHituJbTPJbTUbPMQ94FPEK5tMdU+S1nDQPz/qg4G9X3jabPQOG02ma22raC6Rq0TrXHG3i5q5maN89Km5vWgtEg0X/tQc03mnh75nsv7zFjIAfBc3aKeSEkttbe4FqGjcDdOYWidkrzDVcPeo4VCMllfc+RFkkzxTAghVE97uLVfbiFgrr9YKrTyYe5a6Q2YRCd4c/ftLmomtd2qY+8ZH4/KMymysdVpV2I1PFFzygHENrxRLZLKW7gcVi+zeQWhLoo3Z6zcx3KjGi9vdx96u5Pbf0Zb2t6dGwoNne1jjveUWx2+zkHg1VNsjr4L4uP0TpI3aZjMTcCjNm2CPP3cFjgjZmPLG1wI6ybJJssca96EcFo0cbcKNC+LP5V8Wfyr4g+iEcMznyHqgIRgXZY9WRpzr7pc46o3rRMcWxNyHFMa0BzhrY5ZJhIuOIrdKc6+8MGAAW29bcippJk1l5xGVVFZJo9FVtYj2v78uOSIbjZW5/MobO2t1qkfuGq1AMF6V2DWqD2ikcoOBBzU0hEms4rZlWtHa/3EBdmfGOG0qmC2tHFxNFZZbNdkgFLw3nimyRuvMcMCnwQ7fWd2Vdb/wDaBj1XBm/JEuzJVCMEQdeLq8R3I+2vaA7ZG8J1bLLJj1Sv8NtPqsbLJJTqg4hYfZ8zfFyYdA4UPFSRwPrV+Y3KWCXGatbx6w5JGjrNQF2l3BBzDdkGTlo36svDii9xo0Ykq2Yfs9zVYRtDir8X2e5o7d5UMOkcN1V8LTzXQ0810ajjLdcGg8FJDaTU5h3aapIjrdZqDS2jm4FaSzuo/eNzlcPNzDNh5HSPNGtFSrRaJah0o1It11OjdGCRucugaPNdE31XRN9U2RkbWub3qNstBJJkDuKq8CmQFMjwXsszQB1DX6LH3W2az61plwHyjimyxc6OvVdGxdHGtiNaNsFmvdo4FNfMxvtLuziEytBHTCNuVEHg6pWHu3tp5wa3iU6Z5Htb9bHLwRZIyNrlXm1crZ295wQJcwvPYKdKamm5aSJ12SLGSEbxxCa2Q63a4+8XOwaFpXNpZGbI7Z4oyWUgt7JGKuOlhZ5IVkjL/lKxV4E+Slsr3ezzHo3J1nl3HFpWqdbsnPltFthFYXyHTMHjmmyMN5rsfdLWUc/6BFrpKRt1pHncFFBY6w2eHZp+qq7F3FB8cJl86LW+zau4ucqN+z6nxTJJoW6bOmdE18ZuTx4sfwRbILlojwez3auNAnRxmjP1VwbzrFVhBlc0U1nK66wQ3h1i6q+Ei9V8JD6oNNmiZH1nLRRtDWhXx8FMdYdh3FVGXuYJzB5nj3JlokxkLtlOlY8Na4UuuyK/yF/kL/IX+StLMBp3DduC9tswq8dIzthNkjNWnlqckSxwEWTAeseK0khvVqFpZ8Zn9X+S05mEbhkviI18QxfEMRJnZIHbgmEuq1pqQrmy4YscOqU6zzatqiwcOPfyGGE0gbtu7XcjTUoFabWTe7KvPwAFSn22fBxGq09VqdJJJd4L4j6L4u75KrftQV7N1Pc61+zlGOT7WvNO66oY2P0rDV17inRxuuwTHM9QrDGuJPFcQpdatGBBVOS0zugZsDj3qC+66KlfGSN8Aj/+SmHkqm0yMb2xmV8dO5YTPKjfE854oSR4TR4tKD8jkRwKYfJWiKp2q05A4G49uy4bkLKcI2HnXN660dMCKJ8RtVpF3Cic1rnXeO9HnJytqTzWb111drSaLZcg4NuTRG7I1A62jlWGSa6lS01qr25R2cGtmjOse07kFqjGq/OnFX6PJPBbEq2JV0cq1WPB71oLTsnC8jfrpG4gt396uPBbMO1v9wvOLsmt4lOtFo1rTLie7uVCKgrSxxudC7huXQSLoHroXq4+xyOdxaVWSN7GnZJwQZJlvCBbs+46SQ0a1e2zijf8ph3Djyc43WGTkWOspPBw3r4YrXsN/wA0aWZ8UfE4oTWc07lpIxdY/aZwKDXmrP0V5pqPc9lhP7O3pXjf3JrWigHIXhgEva4qktha7vTQ2y0ZwDlh6LSx6sg4IOdhbIhn2x/VAg4hXZcfmW2FODiC8rRuxschw+QoEYg8l57roRZFqtWeKbZYMnYvPaKzp2nFFrp3xn5G4qgtlpu95XNTT3Rm4q6wl53ucceVtssvxDMx2xwQkZ5t4HlvOOCONGDcgxmNU2N4ed7nMbVHR+148SV/4hZWhG6Jmsbm5xTYoxRo5HRvFWuwXsE5qw9C87+7l4hOAwO8oTOFY2HVZxK0s0UkjNwaF8JKvg5V8FKvgpELU+DR3Tqh3KbRGP2R551vZ70HNNQeRzXYtOaJ0VImbPgnzOwgh1m96M1wvbXJfBhfBBfBhfAAq5HGAOyFpDHce/k9rgNJmHDvHBGQYO2XM4FXRq0ThSrnYBWeLLrlf/qxH8zk4NFS7VXw7F0EawskLvEhO0ligjblfbmi5lmhlBObyvgbL6pjSA0hoqG5ItcKgr2SY4jo3cQuBVpJpuTf0XssZ1f8whBrRQBQXLu0dpYezea/8InU0Ikrj2V0llWs+HyW1GmO4tBXtLOid0g/mg4ZZrClHt3riULPD0z/AKBBoTT3qsc0LGHIPzTZJJInn5ELtoia3g7NYzxnwXTMXTMTb0rbj9Ur2yMVIwkZ2gi6I0a2lwppc8EtwNFgvY4emk39kJoGaa7fvT4ndYJ8LzQhY2pq+Kavimr4kLGUErRH4iLFh4pspm0dw7DghKx4c08jnvNGjEle2zCkY6Fh/XlLHCrSq6YiFx1TRfF/RfFKotJWjtP2g4N7wjcfeunBw3oNc7V/RAg3geSpVB8HEfzlU5TG/wBVzk77hycviHKntkrW9yP7UZXcJAtIzon5UV05ruVW+nILHZukdtO7IQY33Cx7agoyRSSuZwBxCDpLRPeCutdid9KLSt86LuQIW0VN+MpzHioK9gtJr9287wsNZyqTyVV4jnXcdydT2Uk8STRYmBB1q0bYuDRiUA0UHu+2wCsTumjH6pskbrzXYgqrjjwRx1VcbkjM2SKKV++Q5BXPa7Pd+UL4mFfFQppMzdDvICusFB7hbsuGLXDcUbPPq2qPBw49/IQHgO/RUBwV1zxG3tFBotzaDAYL49vov8QHovj0KWovibtUCDW4DlIds717M/4Rx5tx6vcq7loBNde/OnBCASHWBqf5KGxXgKAaQqgtLgF8W9fFvXxb0XstUj91E1t83q1wQaMgncThye0R7B6Rv80Hg3mneobOHEhuJTrNDmdW8Oq1NYzZCjic5zborgukkXSSrWltA8CuYlmfx0hQvyWkO+WqY0SWupNMynenJVuEjcWlFrxSRmDgrU4dremxx4zPwauLzi53Hks99jnYnZWNmnPqvg7T9UeYl0NdjrL4G0fVatllb41XQvVmIFNWiLSKgo2STFh6M/yVlkpvpgr2/cOKM0uMr8+WOd9ndOW4aq1LDLGeJXOWYzHcAsLC9q+FcvhnL4cpriMSKEFNqSbO/WpwWj0ZuyY1Rkd5DinWiXpH/Tk0Zydye1xtq9u14LGDSvXwS+DXwa+FQlZGYy1e2s8JI0Gts9LO44uarxNGrRt+EjOPzpt3L3HRStvNKMfszXs6ruK+Eavhmr4dqaxtkYyRnWaQKrgg0irf0Vdy9hsx/wCY8bgmxsFGt90skaHNO4q9BG2SHjwXRsVWxx+au6GBvg6iLH4ObyAgrm2F0rsBRF7zemfi53vl0NI5voVce2MeK5zQGM5tBRb1dyunkm/GVVxoE03a3DVvFY8lNyElpvXG5UbWqJb7QSd5JQYxk7nHdimyuBdINxOA98hPbG79mOtQ9UoknBXRmg+aN8kI2rgqtSwzN9V8HL6FfBy+hR/ZnRRtzc5NiibdY3d7tShaozSVqo5lZgngHVrie0VRoLnHcE1v/Z7nEZuO9f4cV/hq/wAOTIx9ngFxQZG0N409zRt80WuC9lnBkpsrWja2V7qApzpo9eJ5uHtFOc6EPc41JK+FYvhWL4aNYWSP6INDGt7moyyMDXZDkDNw5DwRA1oHblaLWW1cTdaAtMekfia8krw1hFcFsxrBsawbZ/NNY8R6QYauSF32anemaT2fR77uaJ7+X2iLBw2u9SzUqSSaI2mXFxwA4Dlg0b2s1jtLC1whfGweiNZ4zJ2xkvj4fRa1ticviGJtXXi1xGHIXjbbiFfOrIxy002IGQ9ySFr7l5uqeBRaftKM+SLRMK9oLH7QYV8W0r4oL4gJ0LpQ4PxHinsAq4jBPZePNGl9DSGrY+CpyBwzCDwnMcKgogGjCatKDjbLtdxXxq+NXxi+Kqs78TsHKsT7lnkxBaorILTpGZV3oBquOy910bsDucNyMU1oe0r4py+KcsLU8IGOQyE7RKGNOCc2zvx3t4eCvVvF213qo96hyT54nPuZlg3LpXrpZPVAxukdN8xVUFgqOy4qu73zHK28FpG6R8fcck+gk026p5ZxtPvHBZ8rsaU3cjYWaO63tLVEQZvcgAKu3u/2FGnW4qruR1eKe2J90Ozwqumb+QrpW/kKDpJAIBnq5oNaKD3alayus1nvyC0MWb+keN6puTXNddPFfF08gvjf0Xxv6KgtlfRaSZxfK/ju9wlV3o3tVEsJoMBROgOq8YtchE11WR4V4lYzOHmviHeq+Id+ZfEO9UXCd5p3oNadYncmR8Ai45BF3HkruTWxmqaw4HbHemsdRj1LJWmFAukd6rpHeq6UhYTuPmU0F1BxXTn1Ke9sjnFjDvPLVxACLWaw7SOWiKDZMG7nKrXB3hyWa/xKyd6LJ/5SnCjrvgtiX8q6N/oujcrQxraUIK13gJwgjNO1RSBrsOsKJwuFwB3Kl6h71ga8jH9kqZmgkIDsCGoVYW+IXRPce5q6F35V0J9F0J9EyRjLrmmuSifBFf0grXgrsgul5qSFQb1zkZA4rBw5Lh2XchI6WPEIskZeovg3ei+FPosLNTyXRU8llRGyPBLc2nsogjWCEcmEg38VWquHaHu0IGkGy5OjdZsQvhv0XQU9FlRMDW3jXIFMdK0xFwwqtNG2tduP+YWofEKo98zWVo0m9nFEGGh8VrCnnyGV8WpxDqrBd6pmOCq0+/Qpz4NSThuKLJWFruS11y0rv15McArhfo2cSiY7W9z6ZbltJss7nsZ2a5oMYLrRu9+u5FkfqquxVURaZH3uDE66TTcucLvJf5ivgSCIbyc02OMXWNyHu85I1q5mMuG7cjpTc7mZp7QazuGLjuTRaI5JIwOoETDCYmcFs1XwxK+Dd6L4F3ovaTZtGGnVve5iqudRu5cwzDtPQY4l0p9Aq5FaW7+0T4DuCyXQXvJfCfRfB/Rf4eXeSDY4hGOyE6V0VC3eeQM4qhNTwC1GXG8XK+55l7inBjaCtAmQ9VuC12BQ2WMF9dY1K6AL4cLCyNKLnWFgbvci6OziamGK/wANj9QpnWizsswwAIOapGDKflW6FvdmqurIfmWoN+SbQYqOorVVZWN3Fq3Tt9CrK5jA0mtQ5arIlsQrnAzS7qZLKBOvaHyWNxTxvIo5m5Vu3ncXYqlFPEcsVPFuVC0FVie6M9xWs1so7sCiJGOj8QoJbM+LRlmN7ig6YxEDsq5AWV331rOh8ltMW21YuCksz826zVUbbVeGDm5prz4FbIK1HOYe4rBwk8U1loge09puKB3FaeLCJ/0Kq2YNAG9dO1dM1YygrNAxzCI8UwukbLOBtN3q8DSnFCSKS73BAuZeA6zFg8X97fdvRG5O3I8UWunoR3LpwVtIEPunigJPtFpDcQ1wWjrrNOYV69dNMQrzZBK3vV1/NP8AmVR71+N2imHDejHKSHDiukorjrdIxvcVeitbZTwKvDkqDRUyfw/2FyRte/eF0r1a/wDmu/VY5Kns0jox9V/h30V1n2fie5NlmY103Dc338UQznHfKrmXcFUrVFXcE4mxiQ8XuXwjB4L4cLoQr00QjgG/ig1go0e4LrDI47lrSaJvBixxdxcsBVX5Gi8TqgbgnvgAL+8rRcy0DgquuLqrVLFtRprHOZo83FqDWigHLQuvP7LcSi1o0Ef1WtrHi5GSouhOkeUJXYQx5px0jbg2R3LbatsLCZq6di0jrQ27lgtU0KYzrb1oY4TI+la7lemkujssWDV3J8jXUwUkzj3DxRlPSN1TySUkoG6oXxC+JXxwaqm3aZp6iLhbRBVf4urr7R7WHPrUrAU5O9bVw1UbL13+ajphhy2SsujzWP2iR5r/ABN35kWstBlb2uCx+0nj95Gn2g537y6cqKkpNajlwwxqU01pfCwy9x2mcY2xG9VqN20yV7yiy+bp3hYWmQnxWEjitty2io5b2FcfBHeDiFQ6zpnFGBziL/6qg9y4dpqfC4Z5J9nlGRoqVesLywqt63oPeJA8ZEL2mHFhzRabwBzWriCqkUPELVdp2cH5pslLpO7h7htMbecG0BvVMeTIrFhKqyN7H8VpBkn5jeQEDg4FVs8hZ8pxCuTMuu4jI+9rikgycjHLAa8eK6ErWs94eC5qyvYflCEjQRxaVTkAkcDHx3hV/wBhaq4u0rsPNFzJ4WN3NzWtaGFCkzA3tUQaNZ29x3+9Umg71XcrrsuHFXY8B3cgZdq4+iLm29ra7mhY21fGhfGpssk5MHd1kGtF0Dd7neqnNVebreJV69TvTZNJfDRg0ZEoe0lrKneiWfaMmO5pwWNrf6r4p3qviXeqxtTh5qgtb/zJrWm8TiXHfynicFqtpyUdgtAJdVpxooQBebI7aGKNjEl1xN59F0rvVdI5bZWMjljK9aOIkt717ZK+62PMlCRpqwitU5538vEKOKu1iQo7Nk94vBDTUidId/FOkrVrRWoRJBqVslbDlrRPV6ysc3tVXPQvc7zXw7/qonR83DS9d3oObiDyxh7a4qNrxnl3FMqMacmhc6jiK+CspMemFDi1Y2Bx8l/hzvyrmrMYhTIqn/ZxP7qw+zSP3VhZSPJQOEBFHjcpDXSFp1rvVQIxqi44MZjXv3KCV3OY8MlhlyukOPcmOlaGNlbS6/JEf9lH8qvaAxA7qID2C+aYuDc18Fd/dXQU8l0X0XQfRB0nNmPU1lfax0kjRS9uFVHJdvvoCmODbpIxCx5Q5OncdQCqbbhFon1oe9U0QkcvhqeS6JdAugVRChGbHWM4OLUXNZeG6qYxsWAweTu5cdg+457jRrRUle3Ns1xjyct44roF8OugV4RK62xjxBVXgsdnim6l7uTqCt3MBHV0Td2OKuu2vedptlore4J1os8XMXtWudFsNVWgBXbkXqm6Vmjk7jgVisFiebGdTkpLRZ+eudUJ+mozHVpu962H219/Surrd6DW2p7nHdeRdLJJlgKp/wBn2jpoNk9pvvFzzdA3lGJnRn+JMaXl08usGu6gTXlpjJz5GtlcA4q+Xvc7xWbvVZu9Sqa31QnfGaZhrk6wv6CXWgP8vcqVedyXaVH6lNiikOlJq7u7k2aejAGYhqF6B0jxvIXQH0XQH0Xwx9F8MfRfCk+SdJLAGaQUDU/7PtB52DZPaZu5LxyRdu3clQq3SXnCgV8x3GN1nErSQ8a3U6R1lN53cvhD+VfCH8q+FP5V8GT+6jWw3DTBzmrBhd3BP0rLr5uqRk1SfZ0h/wCWe7lxXFqIuUbXNObsOgcC09yltL+jbUMT7lXRuwc3cvhl8Kvgq+S/w0nyQPs+jdlo0A37Nqv8MVoNpYQ6Z2TuCfY5N2LPDkxULaVxTBSrOt3Ju/BOe7cpbVIOclHoFzbLzDjQlYWeP1Xw0Xqh7RE1n4UbsDKeK6CP1WMTVsgeatULxtNqnWSXbZs94Re44NcXU4prgKSChomE4YcrYR0ceLkI49tjqgJrBoqDiVfnEf7quWe6Tmby1tH5FY3V1Vm1axqBuqnWeTaLaeKnZM/nRRrU9shBaclj7kf2e06jTVxRicNRwulOjfm0q8JBdW21dI1dI1dI1akwao7TLMJm/LuTZ827L2oU4cujd5csf2dEcDrTHu4LQlo0dKUXM00Byqs2raattqq2UBAvtMRA3FFjXXJMqhFsuw461f1QnaOZm/VC8fByunP3WfZ0R1dqZw4cE1jRqgUotLZpDGd7VR1ooVhalcf9oFo702/M2anXGa7k6N29UdsHBw4rSRdBLrNQB1mcOCvMNR7ltjZZiXad951MNpXo426TtcjLbZviIMfxDgo549l309y88+XFYmjRkxGSXGKPE9/cnSybO/8AoqBNDY3yHfdGS/w9xPFzcV8CfyL4A/kX+Hn8iZaJoGxuzDaZclG6srNZjuBQLtWZmrI3geSpVTyObWg3oTFl9jMhuqjO7j6lOb/2e5w3OcqmyL4RfCL4RfCovtEIjY36qiZbosJ4DX8Q4JssZw4cFo2+fLlUI8zdYTRqFnBrI7F5VRDid5XRBdEPVdGPVdGFqxN9U2OWgeMKBNdExt2uJcjwGAQmjwkZiE2QZ7xyUKkLccMFI9+1kFDG00tDho39wqorNF1v0V1twBZsWDmIUdGqh0KF1w0mdVhPCviYVEy0OD5d5CbPH0keKbIN6xyUIB1aptDgBiOKwyTbM3oo9Z6c0YaqwtbWr48L/ER6IGa1CYKrbcGtO5f4iPRY20FfEhNvSh1QQmWmPbi+oRkzYTeT7xxcKpoc69d38jnb9yvu234lOjvXb4u1VD9pGqNftC/3FGPS3fmCxt9V8TVfEL4hdOmvY+pBVnt4FQ2hcE2dkphYTUIPvXh3LDkc/fuRmftvx5NM3poRrd7VozIW96+JXxBXxBXxBXTlXJLU4M8U5jXiWI7xvC0JP4SrxKwVVQ7QTn9c4NCkdL8TIbxJ38jo3jAogzuubiviiviSunK+Jc3wV826+ey9amLhvCmsloku3hqXsgUWHNuCFT5q67PldJm/JreJRklxtEpvPPLpKXZeI3oxylzXDcStsrnXu9UGw2i83suKEjDeYqjpBknWOTBwxiJ3HgrpzCqHUVDqv4cs90Uq8n6+5dOFitR/I/l4v4IuLq96omxN3lCNvqm+zQaXiVd9lY0eK+HC+HaugahLaw2/uaN3KSV7XD0L9WQce9CUHVKru5DrU4r9AmRVwTDZNEyMDrla0ka2o1txrpI10saY10rbm+iDG7uS43o2/Vf8Cb6FVz5KtKuQuaw1xJT7TaXXxHg3vKfabzQQ7rLGdq+IaviGr4hq+JatKbULvBYOT5ZJ74cLrWjl/wCBMce4qoXApsOkpTFCjqSR0kUlpkZR8uI7gjdmuXRdXxa+LXxaw+0CEZf+0XODcbvFO/aNFRf4pIPNf4rJ6oMvF1xtKnkMR6CbLuKxyUJvaoyCaRmN3ci4bRwaE+90pNXFS1NBdOKxtTh5r4x35l8Y78yborSZDwJVX2tzCd15fHP/ADrC1uP7y6d3qoXiU4OG9OBT7Mejfiz+ilOV80De4KaMOydUhYIRjGKLPx5AeCc+aUsfJrUvL4h35lzb7zOKDpJXNkOYqtWR3qtsrbK2itoqWyv127TVJZLnNNLrleCFmjfRxxulYcgjHRR58t6leI4hUZ0btZh7lfkzW9b/AHHtpclpg7FArE62/lv1pRV/yI8gg5uBC+cZ8jopB4HgjHM5zfNdJ9Vt/VbX1WvUjxR0Mtx/eaoTx4sO9Mc0XeKDm8l13qnSONGhCV+EUew3ifd5xgLhkVckg8HAYFdF9Fr2YOHgqQxOiPANwV+P0QmbhXNVO9BYINkNfmW2FL+I+4+KTEnJeyWnpGYV4otjOPHgjXL9eTuTp3b8Am+zXGDi8qhnj8l00a6di6Zi0lrfpJeHD3LjNn9U5pyKNjlOqDq+C7lmq9UI8EZWyiBz8nHgqH7QL18WvjCvjSvjSrrbY4lNaSXv3uPJo27R+nI5qNml6VmHiqFbVE0C1OkdIchuTLLF0ceHiVdFqIHAL4sr4ty+LK+LK+LKMTZjJ3lAGa5Xgo7MwlzYhmd55XNKMEnSR4eKqDQq9fv4pkMTrt1tHqr8GsCc50xqTXNdMfVdOfVY2g/mXxR/Og+CcyOrleqiZ57p8V8V/GmBk959cBfTvHkI6wxBVyTpGYOCaa1wwCrk5tPRX/8AJiy8eSe/s3DVayz/AFWf6pvs55yuGaHtB5ymK/8AtYfzWqECAmPGThVXmYSM1mlaZ+B2AO/entye8VRI2sgqnbdieVk1qjvFpu1XQ/QoGztor1oZe4LViXRro10a2FFLEKFpx7woDZo9kGS+ELQ+OtcnAYhNlaatcqDpHYALHaOJ9x8RbWRutGf5K65tRwKpofouh+i6H6Lofoui+iroQfJCSBmjBGLab0Mck124rBaFh5x6HHkDmoObyXXt1xkU6KVl1wWytlbK14Q4eCdHGzR14NRCulVC7v0TbFGfxFNA3IMkz3H3bsjQ4Kog0kR6wC+HPoq+z18ld9ifXi1PbJG6Jx7QTmOwc00VDyYLIKX8R5brMXIlxqULQahwyA3rHlawZuKjbDM2ztb6rH7QqvjF8asLWSVfnkM0p47vcuM2eUSt22otcKgZOVBsfqroTIq0BzPAK623SEBfFOXxTvVfFO9V8U71XxTvVGclznHK9yF2/cEXOxJ5W2mPMZqhNJR9VR9p2Oq0oy/5smDK8E90z7o8V0x/MumP5l0x/Mum/iXTfxJzmyF7huvLE4L2prtI+LHPf7rbTHmM0Zb105EKSdmO5veULT/nVN5XJTTSYLP6ra+qz+q1nfVYu+q/ZsWEYlDTbXmtkfVXrKwaVgvb/cFpjyO0jIze2vgjHH0pNBRNagpy4VbcNVjBXyXw38K+G/gXNQXX7jdVJ4r7+NF8MPyLCzfwLVh/hXRfRWd7cqU5BmY8/AqGVwwOF5CnQx5e5MJGaRtL12i+C/gCoyylruN1C+y80dUrCyfwBfD0/dXQfRdD9F0P0XQ/RSxRdLHg0HgmMmo6/refBOaYjDcHkjK7ZbkPdqMwm2mNmpLtU3ORvR3yvhz6L4f6L4f6LoPoug+ifEYDR3cuBCFdgpziMdydO/Hh7nyHNVGI5L9wGVqcx8NHN3UXRfRdF9F0X0WtZw790Jr4YzG4Z4UVeSoWnYNfeOUMk8j7tHCoWls0elZvG8L4c+iqICrhsV9aeSzPh4kqqHLJ+IrFEMy48nE8FU+4+T2jQuaaYL495Xxrl8a5UbanuPcr73GSU73bvcuMy3+5dWhhFGb+9FEp7ppC2QGgANF0x/Mum/iXTfxLpv4l038SZMyrmNxrXBURccgr27cPcIKDNJo212kHxdC3Fzic0SNgYNTC52tTHFbX8Sz/AIln/Es/qsXD1VLLg2mYOa591AmRWdt0O13e6Qck6N+LdygcW1gZQkLmqUdjghFJjowthbC2FjGPRYxt9EdGKQVwHctaCp/Cvhh+RTyWSIRkYE3ae46pUtVM9z7rmvQF8eqzU7iLwuFfD18l8L/CF8L9Ai1tmuk9yuyQaR1c6L4T+EL4T+ELCzU8l0H0VQLlx1FthaOIB0rjmo64uAWtmVmsZAtqvkmAVzpkpITZXVaUQbI5Ehlxp3JrPZr2Ga+GXw66BdCuhUbyLrdlyltEs2A2O5aACrDiHIcVmtoLbC21tfRPszjhJlUZFOY8XXNKFIK94XQFdAV0BXQFdCU553qiNmkOPVKMTsHt3cmazC2wrkkguLpUJIzVpRtDIw54zFM0QYqH8K6L6Lovouj+iezRYEUy5DTIY8l4Ko8ws+S484cVmFn7hlsjRf3s4qhhVREtBK0NB5HPrsmiHJJ+Io8jE73X+4PD3D7ruQ/7CPw5D7z/ABUn4f8AYNTfFeXuleam8EFP4+83ln/EPcCk8U7xQ5Jvw/7K0+PI3wRTfDlCb4o+XI333IeAQ8PfCf4BH3T4cgTPFfu++PFFTePvO8OUe6EPclR5Shyf/8QAKxABAAIBAwIFBAMBAQEAAAAAAQARITFBUWFxEIGRofCxwdHxIDDhQFBg/9oACAEBAAE/ITiCW8UoP9MCMoznOM/bPFmCcYT/AFSUyftE/eJ+0T9gn7FP2CfuU/Yp+5T9yn7lP3OfuU/cp+5z9yn7nP3Ofvc/c5+3z9vn7fP2+ft8/b5+3z9vn7fP2+fv8/f5+/z9vn7fP3+fv8/f5+/z9/n7XP3+fv8AP3efvc/e5+/z9zn7/P3efsc/Z5+5z9/n7PP2Ofsc/Y5+wz9hn7HP2OfsM/YZ+wz9hn7DP3GfsM/YZ+wz9hn7DP2GfsM/cZ+wz9hn7DP2GfsM/Y5+wz9jn7HP2Ofuc/c5+5z9zn7nP3+fuc/e5+/z9vn7/P3+ft8/f5+/z9vn7/P3+ft8/b5+3z9vn7fP2+ft8/a5+xz9jn7HP2efs8/dp+xT9in7nP3KfuU/cp+5T9yn7BP2GfsE/aJ+yT9s8Oftk/eP4cYw8SAh+3nv/wBfF/sJUSvCv6q/rr+iv6K8K/qf+Fgf0V/CvE8a8ah/bX/iH8Pf/r/wv/HX9tSpUrwr+yv/AAz+uvCv+Cv+c/gQ8ff/AK+FeL/ZXjUqV41Klf1Mrxr+VSvCvGvGoypX/U/8j/W/8x/XX9nuf1/vqVFx/Kv6KlRJX8K/nUr+mpX99f01/Ov6q8a/pr+T/Zt/0a/yP4e9/wBteF+CXK/5a/urwf7K/wDOP+A/4T+w8fc/r4P9deFQ0m39NeFSv51/Gv8Aya/5K8K/5DwPCv4V/wBvu/1/rrwqV4zr+4/yr+Ff1v8A3Hifzr+6pX/Ef+J7v/TX8K8MeDFeFeFfzr++v/Qr/lr+Vf3V/cf3+7f8LTn/AMiv/Ar/AMOv/F93/rr+V/17/wA68K/rqV/w1/Cv4beFf/K+7/21AV8I8dRJX9lfzf66/pr+D/31K/of7T/rr+vb+Xu/1/m/0agYhlf/AAFf+Kf3n8a/4T+Pv/8AaQ1l3AqDEf8Aprxf5V/Y/wBx/Fh/XX/j6f2n9tz3/wCv9pNPBzTE/lXgf214VK/lU3/oT/mf4PjX8K/8E/8AG92/jX9ARZfhZ/3H+6pX8a/qrxr/AI2H/Mf91f8ANXj79/eJmGBlTj/jZXjX86lfxf8Arf8AwK/668a/4vdv7x4DNX/NX/A/yr+2v4P9tf21/wCXX9B/H3L+4hr4LEO7/wCJX9teFf0P/oV/Tt/1+9SpX9h4GZhFxmOsqV/yv9L/ANleNf8Ax/vX94Q8ME0/4a/66/vr+2v/ADK/4b/oqe9fzr+gmqUS4g/nX9FfwqV/Cv51K/jXg+Ffyrwr+dfwr+B41/41f9lf0VD6r+mpX8hz4GNf9tRP+qv6a/tr+lP+qvGv4H8K/wDBqe9f8Jp4Dn/hr+1/rrxr+Vf3B/Cv41/xH9tSv+c/u96/4RhGRBX/AC1/Ov8AiqV41/BP41/A/nUr+DK/6K/6K8K/v96/4iVjwq/hX9Ff9L/Kv7H+p/5K/pqV/wAb/VX8K/or+HuH8a/vZeAf8df3P/U+ASvCpX/RX/pe4f8AEPgqVMYf+Wv7K/oqV/ZUrxYH/BUrwqV/Gv5V/TX/AI/uH/EQeG3gJ/U/21/TX8n+NSvGv6a8H+df+DX/AD1/ceI9R/xEwm82lZioM/21K/lX96SpX/Ffg/1V/dX8a/8AGr+yp7p/xuMIErH/AKQtTWw847fkEUSFOZREXGDudpZa/NABoXmWCzvJmqjoy1JR2sHhmgt5y/5V/wCy/wAD+j3z+yv5nhdQkblXK3/ylmnDzn22JldwZcromsz/AJaeRAXWPueKE1OAg1W3VZm+R2mAQqbomUckr71MMzDVmH6UQB/3IDWjrEK4QMcruBKP+cPJj0YrV7hPvagdD/USpX8X+Ff91f8AF75/yXLh4Ff8Ff8ARX8K/is9xxmleRuf4U8JFX2Sa1V1TQlyyy8cbTQfI2ln1erFdzbhLQfYnbiF5rRwS8HX6YYKjiDze3h0hgmi8hCJ9SX3sYaNHRmefZzOs9UTcqeSNdl6JyqcM5bhZba93KF9s5mtV3JtiAzn9ptY74gl9kZf9leNf81eFSv+b3z+2v6hALhlj/nr+ShvPduZuDtXBa/rhNNPvCvYKmrdQkcpDtNik5ZqO0mjDrMXWb9bK13S3jQyLsg3a8mkq/xstWerEOr6ELYI4DWz1ePBcNC0Y78IGdiK/THsy56cPRiARyMS3tfqhHOE0G0XQNrtD5P02Yz6bvNQvPpB9FcGcivDrLX+LL2fqRPn0v8AI7K9IP15K3ead53EJ5o62m87VqfTdmJ1exU1c+cBoR7f9Nf9b41PfP8AmCaYIsxY7f8AO03nvtR9t1xR63iEerL8Fm9UNJl9ZfEZQ1fQ1h0j7xuz9dl6JTrrHCu+TNgdZ1lBZmGy9ZrBXdvDoPP9oBjXdd4ptDeKx5l3jQA98kcnd+HMANIilrkDToFS5GtUSoNioKPVLdyIKegqK/Q9Qmi0xtQ1PXrEOhE2NkeEqJHFMPmSsCaPtW3eEW5skdR3jRMqINkjon60AdTZwkvYHDrL1HRcM6a4hChfl/M6G4jifWJq7DrmdcOTMAMHQwYpwVjiQMnk1OT800R3I+olmnj2Zr/zV4V/VX959Z/c/wBB4mxKP7q8VrVnuaxoPkbg/j094lc9CiT9sglD6ARbxStSvfLWXvTgHmAl398EtKxcuCdR6YE3EeI2keIa9j6sdGdZ1nNoM9E6ukuW9R2iJq9NSLpezQjhUBB5Pc/zAIADaWjPSGevBdWLPKDdjlr1Ojp4f7jm8uLv96Zh5TLty7s/Atk/CZZOEsD6vKAAiQMLqB2ZTa8L5bRqdm0Cmt1dujKJF+rv/GNrZNVqS3ugaPeWgbum5M+lbBrNi6sMLo8cTgr45l+cnbQzDLdO05Qd2GQ08x5b0Yr+lJzvpHYeTMp5j3iJgHSZd/Si+n1JWR65QT3zc21RQpHan1n213F9K8kC9OZf/O/yP6K/l7x/Kv4v9VeAy7+0LU94WGqLOGY5rruE940sJkhT1ihPsQuUnPifdKWGYOmIaifIfec3pzAlq0aBK5wi/bjENUuAhrsPVhvyDbf0iW1CdgmzugJtOrTMWwfNJeNwE1Dvp0i8Aluh1H2l/Qq1WrLZa3QNWHjxqbTvPWa7PKGVAeVdVjUrpEpKfHmLjI5YPlSks0ZeXwVfZnzX/PDRLunj3lx0OA8p/qoMAwljtH6+Lv8A5lwxjOOjhgzE6JquIUAJhGahfLv/AIgBojuS9dXyeYpkbX0EIgAdmal9W+jHkqnXWI1h6pPzDPSYXE/eAIN17pDsV8kpcJxOGGG24MQZ8hpNlnmRfT2Gc76S0Kw8mSZrzCdcfRimquU+8L5X6kUaJ6Qbbr0nAD0TqjmUxQ7pT4vTcFxnSyIwPuvwcLW9Ghj2Zr/KpX9T/XX9HvH86/qr+QWwUQf5TLU95OORODc9+CVNA3lXMNXpj7w0EDyA8o8Zt0JsiOsed9IA530Jex9cDlHviB4bsStX0lzJZ9Zucw5qifQwzfSnl1m5a4Kg9R0GCaGBwEfRE/aBW7PqYlXu2AzNn1KQl5g1mEpVoGZz3n3rKBS7RylnSQ8y8HR+Z5e0TJn0dWJYdhp2lzVn5cfmZAPK1WW6xQzs0CoCg7S35UxVsNMvX0Pr4+RTpsfuXFxEaLoe3Lw5zwd9ptmpk67y4/HUNeSWLAvWK8+8yBeJ0894REVjcWmX3j+9NBz1n4hp00SEVabLN4c9/tIXOm5A3BoKJNJ3Jk7kEBjuRegB74L6kvCjiKW+3OPSHEuWyYT3CLzTrNk4OdRJrLHvPy0Sb7O4kDCeoM5mcTbXdRkgZUd0zbnReXMIdTJMjU90257UdqnWrJua7psh3lSzV75TZ94j+TpKL6jPdiE2idmfU1g/cbTTvSIf6HFj/fX9/vH91f0nMylDVnv4mJ16W5Q82aJi+82ln0RnvdQoyLzJwZ1aTdd4m5jreHadWiVrE6oNWMM93zolax+FBlb1lXH6EnEfGU1aXVXFsZOmk4y4yZlMnlXLNdlGg/xkzLluWTFsjvjDdfVRky3cM9GBlYfVsjMB1GWWoacT3w8po4tqi1jgAbpHGr587ErVbdUZYvU9IoxGNMduWVEluVGWekYyK6ITUPurJcsshCcwDs5XQmSBquS3ZZBhHmotCC07u8WvgGpoFwOoB3Z8Qk60fql9GFHmNQwOxf6uX3j1jMzs0e6eesvv6TU39IlQWsK1fZMsKj0ivV5RU4Nka9eqFlp0iP6RGiPKfEZY8IWSZhrxzXqEQLhpfsMz8Es6tqU9yGCY7/8AiViE3EhWPPSfc5vSBW3mitDltMun6wRZHkxjV0nIpnBPDp9ZcoP1Y9ZoC+iN5jl+89zw2SnZXUR9Knc5d1ul6muhaZ7SG02LJhbEh1XsuTsPkidjvmbAx2Y+rUvqPK0w6t5GV8vVPqgMTqS+hgQv3FNbUmteNFHs+NeFf8fuH9Vf0qE9zWOU+m5hl+uJ9YuhGHgmvpIs1JdzI6iHXR6wHJ5VL+ny4jmYQD+YlzPX6KqOINumU4Mcmfb4qXn7hI6G9eBOBeJZTV5Fxqk4rpZ1OoWwvt10QXQ6VDWA4agcumVRDQNO0Qqs9DHrN0BxfeBVi7TGKrQFrNy9hf8AicqNUZYZVAN0jgHoXs5nRD99OJ3eiCrNoEPLdQ/Bl9fRFTw1WDu+g/AQXWNAJ5zcFHYHLLZtcrquWXCSgrZTl0fQxc3L1aHnNPQ8RD6F3FX3lH4Cpmag8E3OhK6eqW4jA+R5+nue8rp6pXT1Tu4XoaMW9H5mg1nl6oCITFLFktZXXz+012fWU8PrPaY7/UraiYRyuGZvXUVlOSAgO2cA/oYHwxHdNljkp/nB3l0OTVNPcTL/AHLRe+y7kRLbrt+coWBXeLWg51MeP6cYihuxJAqA6xJZV3iH+7Qr4M6xtsdx9pueWwY/h2Ax66Hkwx1M+Pzn78IbYpb2K7IaAOXmamPBqWNhecJtz4E2D1GSHUPvNhHRzN2HyRfAjCZLuStPtk+4soM+yMsaHnmcgekVkpa9XA/L6k1F9mfW6Xu8RpJ+ie13Aj/XX8vcP7UE92WNpvg3PVRqiaHXfnp6mP4DiNcrg0FIPoI3HYI6uPVD8QTiP1j+jTYl7Zm1nfCfTAzUq6xsX+BHSi8zK6vp0Ikn67qSiO1Hgxa6PLKYCq8C2cOOfxlcm6NCGCI7RbTV0Y9YaBPGb6zKq+TLLkQ6zZGuOiUzd40gQoqcBGKVegWs3D7Vr8TXC2qyspz9Jc8irTuZkIzQGP5gBQjyjl4arN782Oz7xQNrVy90s/wllvOAMrghW0De0d+WXy9Ep/hLTK1awcsaordHyyzn0xAfZjyV4X3+xLIsjCPN1y8QA523qlk2SPIgdBf1qUjsmnEgUdd7JjiccRgaDDwyQlqi9pZxOOIwyzOi/Al3t6p8Lg1SzmcuyvwuWf6Szl6xFSvnQ4gNcERn/Es5+sf3zUY5m/m+nz2hPLddJiKNC0Wo0Xsh2QeZsiQByR5i3t62X+IZ8Mt70EdB6xvFZoHJK+BzlPrPQqL05mNiJb6469o+aTj6I/QPLJ5TBldZvPqCbDe69oR6a4ndzlUzfR4k9rWSYIGV+8S9APjBlMbHKY9ZR0DyT6COScQeRmwHZmvD1dR0x2ym1DlzcpwagdfOJ9Myfe2cwzXgKZhr+a51O6VOA9QuGBl4Sa4/lBWN3Iy3h+9JiOnGaAnXB+xZn2lVPZUgDv8A07eHuH806moN6rHM3Tc/zdPV/snoBmemaTavJ5iT6FNlGBKExfV3ib4HSHI84n4KlbHfrnIumErN3yy2r7dJ8Uy2r66IsBt7zoTcU+ZgRsW6oR9Fc405cEdDHH5w3Z1jLCGR85sauzPwEEpUVC3ng1nxpHEtzY4dPSAaAnBA3jg1n3k30gWfnM8kesF6Fazcp0Mv8TR5bVZXzl9EAXv0G1mpLzTzZU1bYJ8hBPOaHnz4gBqZB8mYbnpOx6QRVoBt1eCPw8Rjojtek7XpBL8uYHKFkEpMvmdj0nZ9JXzVL4WxTwtAGkzw9JnhGjh/yHrnyh2RJiF3sgvH93xEsc+vYpLi4Vx/tDF9blzc5oRDEvU6S8tlJU+SWggd0fM3h/4PCXEtiMKSeg/o8kJn3t8dXInUS+SUPl32X3lv0N7jqW8vmjjrjtYOV/Q28p34qx2O8OpEhgdR0jmOOo+XiVo+vOzLd2POmmZBnVJ5M9673ZhlW1BKwNHcly+oD6zRuctvqluFTpcPNBoLGbt4l+sMDrwX1S8COSIeaAZu8cD7z2DBEsmLpENnPXJuccfcn0nKQCKuVvLN67TOE9cEOoroZlyHXU3btkP37Ka4Owm/4KBGtO+UcGt4kLlu5NlBynuIzaBZzujtHkJyUdkU9R8B9D8hqwCRixdXNHSPaEqmjT0Zr/B+omqIeCI0FrpuL0p1amip1XNBugHgjtRDrFe92gaQ7oL/AETU1kTYktlIrnsFU1z54GArxGhJLavthBF69VnPeiub26pW1XZVFr35W5rflGb17upuA6YxCzXlbmzvS5ybyCbhOmMbodzlh10urHB6voes4v8AhmJ2O51glrUV16AesPUpZ9Zse+qJDvqLZu/XL9U5B5as7kZpKaXKzZnjMv8AEC03dZXznYzzdqHltXpG0IyW1eV5y+L6RNhNVi+xuazs+8pqW6K+4yv0xp/mXgQ0p+xigysTJ1nV+k630nQ2xgcukW3kosqdd6TqfSLbnVDLaEv7CxdXjsS/0S+X0lGB2a2l3BrZpsekPgRZ0RQMV8oy+ogtbD83L6vSX1ekXq9JTIZ3opc31xlaBsTvn3Hv4fN4HWXRPKfeBZTsZmczm7X4T0YJEZb1Uti1i0Eu9WwkHadHk/EtFptrMz1ZA0rkYuE6AbfO8WgE0Rnwsr2604Lyn0OZbGPJeTuS+D1hIhajNefJ48nafUeTtzB4EpUR2Yv+BPlBnkj6u0olRuMXgiju1xa3lK9EPhiFkD3lPZQl5mqg6x0UHexSCzdFcPO0z7vh6z6KX0IVx/SPXZ5MM5OcFw0g9coxQXBwwdDypqW6XCboXkYV12lTMn2mOt7U2XflT3IhZMCdNUddX5xm1RL6lSJjs6o5pXfGfTQXDdq6YmPvOE569JY/MR+sJUo1fLMXTDpRE+h5ELLtbNFHRX4Lj1pXP3sGpBGzcSvvKwWre8J/CbIXwEz1vcqHF8tyr/km7Tul3t8bCiN5fQVDOt3ZhhnAuOvjrjK1KdDA9Wc5Sh9hEv3BwTcgdMyz3pAGKvKXqc4zjpgcq5bX6Zgh+iJxl4uV/W4pvg8iabnzdsp21OqQFTXp9ZtBxK2OWvqKfIzDDsNs9Vhz6SxsdUx6RIoqcDEN0HVi2yuqvVNXg5KJgGOk+NmTFmmVeUvSOEbf4lpTbqm1850XrLIQNVZYi5CvLzPX89OxtOi9Z0XrDYN2drM52pWPfmFDADvL4vWXleyrRHVO5avtjrC0F4GfsJ0fVN/s9o5cEXnJM5X4nyMvh65QnFqukqCLkcfnOyL4RcKHcsWx19dISAAYlwuGFQFZYtWp5rlw74vl6JnkwdOBO70T5CP6kKpUuDQZIBcS93hlf5oEaIIqXYNPhZZt9JfH6TsQ4CDqqo5kqKeymVwz4CV+qa1jUTVck0+iqx0cGA/8ws0+kcsg7VHWzq1D7GKLsCuXqQP0x/WgootMT58wRZ0e0NoKrRokty9J5CxIiynuZ8vynSlzXk58oA0pZ3xR3O3u8by7v66pg8dJ35l700OE84/f/wDrLYeheukNQSXJrwwKXoo36I6o5nPpKsKvQHlPmZYF8hTDbP45J9I32JdqPJBNetH29yPecod6SzXBsYB7jvFrL5qpvo8R9crJh9fJph+B5p7YMj3lbh97T3fantDIBbJnzRLb7pnNu/PvK9b6MSe/cq9tvNn3WJXXHVXDB7LGGVTyEr+4uP8AhpNx+6aG/nOiesAMa+ulbRgGqIFmC4fnuWYLpe7bm7nZqArzcrAw1cDNzd1UrXT4jlYhwJ3lboW809wEt6vRUQNLeblw1kOo+zSPQ+mWG/P1wQwRMYrcGWD8PIVP8IIeivO8Qihw8RuV9A65Qytd79oVUAjWIHWXq9k9UEYPl5mstzv4RFxtn9l9ogewjygEoodp3Qhi2htj7tQ/xCWouqyvnK5npFP4I8EHUHrMOg1CteRv5wEoQdp3npLMz1WNlDz92QmvsjfcZXF6Tsek3JMAWnATAQNnp359oGYHpK/XH5krj0FMH6E3jWTP+J8ZPjI/Mjy3MPy9YgBQOk+MnzkwjC1iIt1Y6H7tZ1M6qdZD+hneVS+EH4ojqZkJn20vzlpKkqtcN2zF+d9blvAC0kcVdC6TKKfampLw7k7nrLqB2Dh1Irstg6x/ancecPNNSmAHhpHPR0dYAWMR8jO/1QsbMnPZ5JljMG/oeky/JEO76xJSqd4wtt37Dbyny5ktvDrR3vWFq4yW6TXN2N7bvOPrA1xCfC58biIjLGT2xPlvLzR64h5T43AkAOzFrV8Dfon3Ev5SycwXknagVd5nBTtvzOfHyN5UD9HwSluZ7T0njPqQ1N2PcJSA8xSkZwxJtd5XtK0ycZJv3rS/UQGxeogdEdSbl6Rs9GHD+mU3F2MesM9CZq8ed5vzowTeD6qYKoX6IVhejcSuuRhPxpubB+ZWqzdNQwQ3zmW8nXU2m9Bc96DhyV2JS2/WdNBup63WL63tIuwO9yxfrKm1jv0vFx94HEo9HpmD64AETnHi5zTrjHVj4MM7AuXcRaGXabeDWbYrnGCsY4M3g5ZRSC6t8GWbFOx7Tizsp9nU6vogOleBbL/u59IZFziq9EOxEI7B2mlPWzPpvXDPceXtKNE9J2fSeupEIDYfg/xilHpNxXH6Ts+kOlwrDDSnBe5gFUtq1lnwkx/zLUm0O3z4n2hnzby0QOlCfASv1SpVojnz4IbMsi/ZAdKeU6z0ic3pLEu3XXgTTzdnkjaddOunVzy/7R9CX4Pbar8eKczG3dEfUcKT3N13X+FWGCL1Nh8EA7KgIP8A3l/9Zevuy6Gx17C4QfEz5mfAzLDOuj5GfAz5GfIzDQjPvr900fcnd6pXn1QeX1lZIfXxtebSGOr6wvu+sQzb6x3xE5mcLMwv5KHRad51H1lXd9YvNcpHdyz5ryv5PomGbWI6yhz6w+TC4LqpdvtLv8KE10gZ04XrS3VncmW0dfTakh0Tc6JOmTokvzDTQnZmyVbsH8wBw2lXcJwCHGmmNNMQ859tCeejPO7GHQTpnpG6LbiHnD2pr1yp6FKvs6MOAnTI7Y93T0JGn1IKEnJ+rSMrSHclSwh5e09Jwz6k0HTJ7hKcjlSuUNdwtpsp4L95vEdj+Z6O15lveHcOQUzY44b95zc5YdoLsGWbkz1JyqZ9g5TZ7z9hjewmMC4TzmWrkKpf6SW0aQLSX0wf0BmQoPJjwzb+V+cOA/xLHbjvbN06GB4ZKF+YYt1JOk7ttm8OjAn0/R1wecy1Y4zlfHV3Tf3QNPAch+SAqbcBtlrQ/BUS9c0lT0SX/onpBXLvqqk1Np20p12HwnuK6vhtFuyexesxBPTwgLUk+iL3djXRngrP0NZ3x3+iHZd9P+TD89K7/hM4Hq1llf5J8hLKBdC3YJQbu8ElSb9WrXu+CKmLrEwQxf1PH3Y+K6grTqzo46P0iDU+kYsDT+i5YTGtQ2vWdN4Mr9Eqz2/gfQmc00mV+J85PnJ8ZFetYEzsBGbHPj2jPmJ8xPjIFqoatRs9mhs382dV6TqvSdd6Ef8AAIC2Sm8ar/J8onxSfDJ8EicHvUYOo2jaN/8AWPKKO5lKEx6p87PhZ87FCCrXSXND2W3mljOTrKv5J8DLmDUreNSDI06/tP3E7n1nc+sdYoOyxGT8qz8GkoEiwRTmFOfUmre5LGpll5vD1hp621n5Os+RTueqAP2xzy469+SVeRwt5kXQyO9pfs+qdF9UYqvVQ+cJzj0T5b+UrpRrb1CdP3nTlQBte0PWgZ8vylIlOy9nRg+yHEiABwSvwEePxPp1+1qSx3gDDUodpjt5cT00nrK/S6Stx1UnB6UZpL4wcZJ9Z7ej8TR/ECyWh5WU6D0mpdzWZto4K/mXMPI37M7CFW95fsSsG9Se2YbPRnCL1w9VeD1IbY/RjjoTqR1TflVNtHH3Cb/7wXqvYX3lPiM3UeTDHTDpin7X+ZjFaJg1h1Air8Ex5wBcU0J2ZsB0ojOs5ymJ9qDXh3li9+qibkp0LYazMg0EdCNNZVAcdtm5vkYl/SZggNP2HgWJUdYW4wbVflmZZepll4KN8F59CGrPkQS62dsubp1nrMXesJTyDn/ZBFjddemIFEbCTr/WI/6nVTTad+J96K8/wlch6M+ZnzMN6TqwqV74fDeLb01tL8T4GdD6x4vrGz7/ADi2h9BZF9nfuwPb6zoY6H1mCcW6CaOd69F04IOOIAz9tP2U/aTcdG4P0I55z2X4l8fVOj6p0fVKYplVhGARG+HaDC+MdGOjD9LXWpuekFdAHiTcaMPerL0wnfGrX0Tv9E7vRKm83NT9JPkJ8hL4vSI0ETiIYioK35J2/Sdv0nZ9JXH6RE7rU8x5RBMrEJR2RVZcN5Mwe0SydY2wW3Piyv0Q/Uj+pP0csUZdOOrql3N1xkeGfIT4CdV6QVZ3wI6h7QqXTgwJA06S3+ER3y1a2oBmXb1P1SKWhqFPlzL5oCnFxid6G00pfclrP9zN3lLL+g5J+zn7OPL01MiUMYbv+pC8UdVrz/MACRuRrmerFdUPeVa9Yn+zpR1/zZ5xOU6fUg8+qVccGUoWp3vZZuLkL9tZb5dyaTylOX1huXFVPmC9pt/sD6krh8cZJ3Ciydz1lAI4ynsZR9DK8w3tDL/YWMyY2dGXNVHbHsj6k3SnBHFvJftFLeZEGLq5QieEiebHyxNovBp9SW9RYp0/Vl6GB0o1la6XTKHuBYhlAOkvlMSF8Ms37UHEzsRWwPcMsjySpPMqetks+k1PSLog1E9J1iH2gOrPo4X1gfqY9Ux51S2dUnVJQH9WfAmesPLv6FVOITpvWPE9ZvqaZl5TbF9f0zz61fqdL6z9lH/al+HuXq7S5YL1Xn+HhqR0XrOi9YBaXnBJiwrXn7+UGFHS/aj99OnnRwwt3UWVuMPQbd5VEDld1yu86PxK1N3ArXgJgI87Z15sA0fadb2nU9o8r6QH8oQ4mQIOUX4nd9J3fSd30Yjz6pTAY0dNu9iMhUAsT5lPiU6XqQZp6kEQt6eb1nR9adD1p+5SkSEpf0ILNGV3Nys1ZKwVYKOkwi8fT8ar4SfCTAU3B1ifCT5TwFpUYxUjvEvbEb8PKX8Qif0EoFMXhcnmsHDXQ6T4BEP8o9wk8pduiNu9OL7PWMzboa9Z1/qTq/UnX+pMeEpVZgqndw7/AO0xFNEvK4Sbl9SA3epPkYCsJoUTow0q/wDTN4ZZu5HSx08P7ksQ6afPmUqL0X4bQBV+9s6P1h/oS2FB2WMvRJtfHExyrfb5pqSrWN7J+4n7Sdtgyi2+tT+clum5P9ccm3eyJxXrmKT1gabjzlvF8xumlfoPfPvGPmxXMk5xR/NavaHb4Cn1PxD2mvdJ3c7LwgqtOpAu25XXtpKuA6JfWOPUQeshlK/wRBQPhtHUQ9HppMag7ie+L6wh3TwI0+k6D0mn9frxJkCBaekbm27nJ9J7CDCHZLkJ08GyAl/sI3Ng/ObB9pOHB6Q2j+BU6KakEL2zbm36nDKLlz9tIJQBwEOHM5D1sa94alwH3dJQIjHSek6b0lOyNH8Xdd3afWLPNF5YOupd2dAnQSrYlj/EXXd2mv6u/X8J0aSJXiU4iOJcb3FO/EFUeprzN4JOsAUEpERCWpL/AKlsQ8Atn7Ru9WBUqUeHloFuvAj103YcCV/DhCy+r0m9TG36HB/Blrrd9z2IDyG7q+rKleN29NdXfymkJR3efHHg+yg+bUEfQ/Z/CoPgGZ1SD/EaMan42jSWc+NSoInqvnzTDdXJw7kwaWypkphhtejOkrE3gBsDddJrk27cXgx4YY4jHjaQT720dTklkxCITStbTyRvMXjqfOUCVTEQawWxsi9u7/ukIIuMjz9vOCLGxmJiUcxox9dHsaMPqgfMakzpSFSvJDkJ1iIVpu1fc0Zscv2vxnX7y8ncnUJ0k65Hjuoj32fOG2v9NozCK64jyYf7k4H1j/rT4whaaz0ovrzESFW2wHs6QKxDoz9lP20ruvmomD02eh+IY/Wn1SB2LC/80s/JMI869wjod4r9ybCOav59pqierPpDhzp4t2Uw+s/FD/M/SwCjBDkuYPmx5fpA6C6PhBdhOWNGPW/eUzF3uyGZl8r0lCgujP28q1HzhVO4lETxKw+hB+X5B6JQE8E6PqZ0fUwvya1zvJSntDK7f9GGQTbxa0EtVYrRXy3L1r5r5nMN8cCdb3Tre6IP9Ir6O1ru7Rru6bC+8V4rtD9DK/wxP8EPB+43aJoEu1i6u0Tqs3PefEfmfG/mPyP3mtzz/RBVn76dlt3l5LMpZOVnRx0MdDCO2HbpX7iYuWS7N+s6fx3DK2rkerq8E8hxl9A8arrPSdZ6EY+S3BBLFSHyWfoifGJ8wnxCfp8buWeMrVD+F3dqmJG9Gha+5Lf7y3+8+VnyselgtrN4nc6T4WfKx/dh+/EeQpzFEoQ82AzVnp4eavyYBs1tfHmUNTzSp+6n7xP3iPN6kM7RSP8ASbZYr2PDPmUP2k6XqR4PUlBrlbZ+SIYl0bV8/hDjfWdJ9Z0ffw2Orqcj0i890feHWU8lYmHwPRzpokb9QsjZzVUx5tpT3dBSduYcTwLoon8Ewv54+8N1PQvLvARr0d0/TwjrJsMT0xHnH1pwP7Mp4D1pPlLYVbfSdP6Rr1IJrSTsU8nUiwp9Hwd4j2beP1k6b0lUAdkjLg77zE2OP0L+Zc1cX7DAO0B0TPZPPXtvaMeRk+iBh2H75OqHFcs2lOCeoumfWfBmdcx0hyX2ZidwPsMG9h8Hw3MvBnqxwepij1Y+mTNLHcSuUCjB0lJgmOLoZfSH0pHtrMzC+oEdEuXDFAOWJvKX3NJhWPe9WNXd33qmKlkxL7c6G72J+Ub5flBnK+l20QBRgi1LiIsyjX3TQSzfVKvNqYLAdhLlkpE4Bupo1fpL4axRN1T9V4qeCyNdPcLYhUxyPtG71YJLizGGTS1NIubqaPtjrB/BQQMuXEwTp+3XV4Jjxqrbo4Ig3gu87pXmCbkeTXyJ/YlCrIg3gK1JXkgG5D2s1u9JYIadQas6hKNkOJOi9YF96JmqjMD/AH5+7jbXhlP+QhlRcAJSqcg9EP8ABz9Xl7XsZ+nx/wAjNCoGKNKIL9jP1SP+Ol79pP1KMhVmpewyyCM5ym8tPlCGGg6iZr2U0b0kx/bRtjQtrpfWAxQ8iH+cn6pNePyQQ+ylXMNmW8jGJ5tvnOGURfJBcbyVaXljWKHbHgG2IffIvG0VZSp04A8Cfu4NYNBgIa4fTdGGofB6Cb9yGCF+QiaNmoDL9Pm7T4fxQt/UXf0ilsy2u9T6T6FEGDUp7m6UPtLOeZ32nz37Rpv4/acGCK9AxMGB+HV+s3ocxHoTfnto+kNWPcz6TF8n0l/bnz2gCI7JfWlTSTSxeaPpPm/2iMM1ISD27Rp/SfPvtEfUprEtmfEWT1i3Xt0Xrklvyku7+3CETFok4Y1T43S9p5paXo/EKO5IEZQLZE1ukMaxDc/1OhBCYNQf1eanxH8ylkDhsW1NZwge5ma4AEITRHWTjioXG6V1xHaFaxfMCkLpFPvC8p1J62rLYHcHUZALVQjDa/3ZBh95Xo8HLWPIiOMRy101QJt7kmgEdQZx9oe8R4vypMRUr5/aXXVnsbFz8DOKAY85S+P6RKH7j8ZnD2aN7TLs5pw7qRK86h9AQk6RfPsEc6gHcMUTB8r0joD7z2hQKOAr6YmRU2x5lZmi0Qn6IU2av2WIg03ejyIh+L+JwQym+wqKBNa0HVV7ShN9XomIZkCwyXriYC6X758Td22G8285fXRR1orOkPQndQ6vMW1atgXtBwEG0sGYfORj5lRF6HrE4HEBla+DMZ9HVOB1YccWKx7x+C/WWAxpnpy5lE93Wl9MwW/z9Z+87TkMZ7WwHCFSPYT6yv4/vH2b5b70HwYLyvrPiX3iG6upc6zC2ruRG+T6xp0+r8wMdas27+IAiXzT/UsMpkK92BTdzOU/ysf8SGuqoYvfgKpM431BVK0gAdgeQ+DDs+kiDYL8S/kQ/wAfKWPRzFa0qx+MFaQwton8OKMehiyqrMFqfiFf2M/xmGPx/oOGAGmmXP8Ax2KZhThG7qpbfi4o+2gtPSSyyy9+4TV7Nj90/wAdjfg00BjQ3mwIktEGYnFRwiI/cT3p6JsZ2sfgfA5GzYFK5GHhZp59EgGCwCmF7Gk1S7Nsr0OSIB0atJ14YQEBHclUC5Yr8jKtZaYV0bxCd3jX7Qdx/itXzXA79mbDupovrxEFQmiSlRqd6iMU4dN+5AW5Aa9xHXAh0m5UF9ezv5wQa4WpRaZ0SyYLPU0/mY2q2KL3PKW5U1WO4Ti/1MnZjNf5Q/maAcaUo1uBz6TtB098gntrG89GHui2/lzK5LkZOzGfW9dA3BDZMhRsc+ktf536WsPKqxTvowaTf8R0ZqJeOfWLesu2CKz6aDAt6iVStu+8TydNXoSmCHI90lzNeJfrGe/WGhANXt9JbnPK8/Qod2+sveKcC/TCOPe7n+nhakVQDuFe8Wrlg+qPudvqnnpW0F7sr9EcVTp9CgHqAlSR+Fe8veFGz10jr+/uZ3Qi9xjys7LmONNtFgF7rZRCJDxlpXif0TbC/udCLLc9cr5zvVpyzQj5Rg+xAevmF5mAg/ZqHP1xRNiWbuTiyG6x9VBCDVKJs/ES3oQpTuTI83bygV7swy83Ws0KjUcPsd4751fNstF1GdIJV1WtunLA2cgnB9k2ESEDia1KCUOlpMPuneRNaFbL6ake0MYLjqhQsml4Xo7Tbmgb9WKEUX3GxTUgHXvbpCHyoIdDTm57Iigbi9n1Q4God1yxEI1pnmus6hSDsIT6IEJoTIuptHe+45GMU2EQptF0wccmxKpWt3i1CNWBdFhMjMthoA81mG7LQ3xDvTGP1QWsHKFc9jQhV94YtV7wrfaWZwcVnT7QEmkFY7z25DA2Ayw2nop9WIzA2uM2Mm2GWGnMdWCkpPEcqxw/umY85IE72AMK9RF3cxtvgtEHy1As6yrJXyoJuegQ+dTWk8Vj+1rDKM1JSOg1moj1MTTdB/oloYUMS32l3ZOamBX/AC1ig2DENHMkEd6iZhoVK7+kuJKal+JlIPKuBIKvR59IUcdgnWFljuO1gnnKkXYdKPthUrqDu5FgNCx9F+UEaq9g7QKwKDD6kVVK3D1J3POIHlANDOMntG+dpPOVGvrYOyP4plFnR6zZ8s01Tz9ezaH43B5kMsL9YSqjae8yI+JyAs7XiHo7YPc3gtZ3+xZ0oWF7Kpjo75WuzaCvk8ItgG8dmH2HVsPebTzOP77k0e6IeW6hEI2U+eqYsni19dhmJ++RCq8bPtY2HuSj5VRJhUmz+8oBDV0PpM9MaNnuM/QxxJkm9bQl85d02Vp7Rbrsap2aJZ0LkinyuDZArsvMmSo4SfZAcp0KL6n2iCjbb6omHS4IntG22v8ASNQB0dUek5eer7MolUznPpKWwbP0WoTYr54kuCGqbXvMNd0Vnq14CFRsGca8RQPyo/VLnBJLfoYK3Op5htL0CyqQ9aRfwi3qpgOX37sCpZ4wIvsiKZ6FqetyvR8/7ELW3laum6PCuXeykrQgYTemYQHW4PlQRk26NL3WWIgJrYRCAWACHoYNdDoO4oJbBrnbd7jhozUfutxnZcCC3bVKwRFDR0HSVBE1sRu/KgPSPQP4VRRkDSdoiie2ieu0UbM4/IpC97XmXzUFiGortR57NP2jT76+5KLi5X+QTYfSCnQfxFqZZxD0CNDOjZ7XmFb1n34TakqlYho+UYYktOKTXAJmOoS3p30PaVaPQSfYRqav3VGHPtwMDqxVv7K9IrdbzR9ImfibmZprRtXGmWDQHKpPogizR8i5pYAy+wwzxVTR9CWtpqCuJa1fW+mbfwuGwFx1h7YAvMW+DXWC4jGNrYi7WvQXhXSDQPal+U1qeWJD5GawmIWkHiXLmHUCz6yhiPNbiZ2i3VOxMVTywKxPRcTtF5o+kc+uoO3pcZERSHoGPWO8m3vDEheFREWqepCSqNxb1nt7rCa8yfojxfJLAn0Dfug1dnCNmIejW0RUbou+VMF3wmsR5rMkcGVW1if+iOHWE0P2IMVMZQvvTkAA8bQP3MhWX2rAVdS33JsbbDcArSJmP38Je76C/wAhUobWok92MS63vNBiCHPQcPECaEKEKlbkSpynL5/aOqfrB1RF6SuGCVquDzhHpOT0UxqldPBHWdDX/E2oMtQXVNUanaULtSzbQr6fum1KS0kKgMAmo7ykAM8XtBy6oX7JpkcTMWcsFY5uCQul6A31mkyZLPBYE23EemzbrHc3mKgxfV+JQI9rQGKjlZriANoj8EYJFBNRiQtwLC9SAUE9AfUhMS9B/wBlEv5UkM04hQ7aRdUXReihKznkZPOVy3IlejBjbFyn13mbGKAW/maq/cfN9p80A1NSdiQMAVAV8+MxPGbqfSUPl4ejL0KzZX5mYHYr9Y+8E8VtD20QwoDuRG38ojHV37JPODmjs/aXukFj6GZpbPvVz5z8yj4qLaNZSvczF0fbVsRS56T6S/R1eyh/gGqKtWdqR7Qa0X8JtM00M2vrpLotlOSafad9ZDGd3fftAwg0Aj8xbqFvy6frEcGfGO7L+baaS6c8IX6EBM2QufTaHTcOZecCIiHdTHWe3XkNWWsDnU8htHB7Y3fKcXKrXv0gW55y900WgBRKqKiXSf0UVGv81ehA+1TqKuAa3nEmZ5DA78wyeeP0hiLGHM31X2mQm2/IO0uZYbXMadLGY5KnxToQKg33RcKsa1do9gsHPRJ+/XPVlM11tgiWf8EIwtoluuDp1grQ1oDwBMO1Yyft4c4wzF9tBzMlRMTeKBm9Oj7phLqJq/r627z1iCWE2oHWWBuzjHXqwdWkKNDILbtBlwUGf8yAANJWmt1Uf+zuMa+cvda9Aym81Dn0lxg+cb/zwNuSlUL6drFmnMshFVNlxeupMehliQeTZdvPe8S5TTcqojqeedmYui/031I3Q9+9GU6pcQXQbwmtmHhaDOqajNJBtpbiJ3BrBmpFgfvnTJKwP5Z9oBSwsfAAkKViHNs0f6S0FYew+8v1BuxeB9uI6dSL9fT6QFyRYwA33m6TJabEWOaYWpnhTiU4fYuPXSFv1Gz2eSBCbL6g+BTePBLnek1jsWyNB7M1oIxFeCEVqjL5ksi5pm6/yJXidd/u3lQBq1G07ONl6hGxJx06DAusePbwRaIWuO8y6lXozlPw5i8jwjT5cy4LrnK5x47UvUSrnTPaum8XS5sW6OjAEk6vnZTJkM40+8th3ATsY9cahKmqAtSnppAig8l9YukWDL0gi+bhft+J5iA9h1l6UNQhWboI4x3oMJt77QWQ6/gRYYXZe9yVc4pebGMUfH+x5T4t03leY77Pp/tcYD+Z+ufmYYDkMHUoTfNjSGky3ftR+IYhvyN/aUs8TfUS6gdxIehcfJqv90eqpRXOPylyrazO2/QnmYIe2kZeK9d6JsV4vsaYzSvH2CMUchh5BLkW8D2FnvLHTYB5GrMnvyc9BjRO3t+VaS0FddD34Z7JyfT8pcpECroXjHkEZ2kRXboSloR0z7+8JJpcR5pyIIW+XE3asuPpM9Rhew2TmsFj1DEYPLiHGw84NftT6jX5gfV9De+vvKvraSDpnWdar4stOay/Q3Nl0Q/cIFJOtXrDEMD6PjoTr2oPzR+ZsQXUe9fmDVkP6ic+Q0eU1j/bPTSe9U3qfiaFBGkmsDdNuhTggn1oMHlgidG4/wAkNOCwTslRAZJZ0kWv8o+mOjetfcqC/WwfvFIXdh1MwMHSKNH0JY1AUegolhBw15p9FCDmYZd7+021dB9cMIFX2ISOWavkXznoBe5P4ij5vZ6aQK8PlC7ssOLXupTF+cSbQfmXn3gjYUu12YrMaGsHE+o9/V+J1IyP8yl16lBn9QBY2Cx0mpry5es9yT2TACIXqX3hylOEZrNijp/dlunJn7x7wngNHmXd2DWdjKqNOSPpyv8AQxdoWjt9JgDG1p6IczYx031yzDvvf3ghN3vNJfOIOiMjXhNWr5fo4iqJKqvmRyslZXuEG8qKfmdsHr9TM8BBNiZx6BmOQ9C+h5S/PVH9mkvC8fcEbl4vW4CF/JTbMco+cv1QWlWOpEMKYG+FYX6Qv9ICb6M76Q0DQDo82VNP7arxzDK6Q9kTU15DPrAqCabUHuIrtbW29oMWNy91qWZqtNrkcMCiL718TLHI0PyiieQHhKgp0IYDfVsekOqtGuvRlWidsjXR194khsBecvBm/wBIlMN2JSMD0UYh5xCMZ5B1jtTQMFfcie5k9YLMYq+udc8O+6OhmBUoR2nbG5rUR9oxyoNPuIABTDT802+Siv2g4wkto9nE6eIEConA6jZNfA7+xB+uymvtNpmgwHoMMsegh1m1MV0PZYhjTg8AGksdokpXrobgmur6Os7gltXmtIaRhbxdfyRKwtLF7QR5VfhjT5MeUHEXTKQV379Rqm2X9jYgV4K/M3hhe92xPRZQCBGIy+Hmy59JZJ2p8prUW00dA46zAmDIFlqjbgOVPdTRpjDkZ1VRHXQ10+ZLYzXH/mSlmDSPOasTFQECteRuxDMEWKPEfMzScyYzenPeVlJz/SLltVWU6wGpq0wd3eDwBoMRiygFxc9S1FcnKDgdlAjtnp+CX6VvUdkHGGruuWaRYAI9DdeCKeKxaet6QpJ0CgjBQLU92aQXDt0IboX8MhBhBhWrtL7W44IYShKC3RLnNcT8CV+f4HfxK9MEDeURCbUS26Q/61nLux0Q/jUrHxbX6sNAzLeqVGO1iedr7QAFB53hRBc0L2jGOini6sr2jGC2/vmVKgiS6hrFb1h/EG+13t4VAMtM75IESAYARwfOeJbLHqt4yNoLdEob/CKJYh4MF75L9QmM4TrMDIfYJqQKzQLV6S83stXrDwEcOk3lEFV8PSLbCwj81BGB2dZXhOjq8ktaGE0HDASyV4IZgfB6x2t6tIwmABkde07NGwlq1OPMqAitqb93i2MJO3aZOOUfNmfeneFWUUkA0rUt5BWIMfUUGzmVEszwm1h7kuxzFsQtRKplYv7VByOrACPWLXRDbBw6eFXESds3F913pvJga/sRdcjBFZjZQ2b5hK8azqBIPJzBvwEl7UvTY4IuWjtNYord+C5d11XsbRC4mTb+8I8mq4SrnTotkecG+NYEWTwdtoYDdTo8/AEYlKGg2lBGqlDzzBoR6n5i1qaUPmfeVuDLD0FHFRp4JxbOqwARNzWLv6kLltRMsS7U8o1Ielk8zT0gbM7lr5zGiN4kOdUqLnrsRhM1/S+sYQuRYp7y3kYDVu/VM94xSvT7zbSBWI0lyk60byokjksiAnEKAdyBe46TttMk4tWPWaCGh9Dhp70SyMG3BakIUxPb0fmGN/kDwECcW6E4ylegOtgcrFizG+rvC6lwU9gxAoW3VxpLB6YNVAukJQdYyWE4p9XyjAqKf5Slvgb0glSNU4DBoXNmh7aIXSEdyEG8HMwDNg0/UF4J1jzWswEW3N5fyitMXjXiVFO0JqvBNORSxeejAfRfby5iMjMyiecRlmXLZCXifuu7oTe1IA2LfaB00B9T5wqkseggrH/02jO/WP2GMOg1J7v8luEtVUs/J1ee/lH+mB5b33YSOorW75RWO2kFbsiZmHPzDz/CY4E6vA8pauh7QlHwJpiLQ5XlNsfLH5RK3BYK16IWEfL/ACKAksjWmO3E0z9tfdOr1U5JhGtp2aYVzhLifoL93E+ASb6Ep6llhdssOgFuD73d36iYX4g9yYidFXmJXSDeNyMDPVVTPX/Bf4jkOfvzqzTRem6XdEFaaPeUO9nCHjce8C7W7snk+8qiJ4Ccy5MeTh4nYGF18pgbf9LVHNH2x2jNZbDz4gSr+4HzIZFrsw8n3iv3pDu0J5X1qcMOwcTK3hIeeQ/SJQylKvycR2821nQzkACQSx7n3YdLl4Q1OvQ7eZGIYmNfbmLQAN2WPC4w76Itsl6/mUDe6t1+bjqXgGfMS9SNva8xxK7Xr2638pvEAVFAwh3XuE78mT5wV1uz5/FtvBrfRahhFGK8hJajuH6ygl5q6f3HlKADGKn0NSEWjRLmNNWmU8iYJz1/L+UHhNF2HbRMaXfUJGxsw61C4xV6eUSQLXNvyQTYrTlAUuVxFQNjDu6E3Sf3G0Yi7rlfNixS27gFjLolxDvGOjzIUq82O8CekzBV7YEJPywW+01JT/QdWdqXErwjhNyEPpChsAD/AGLKSWvdVO5oxuiP1mjGmLqGeJROgvYQzdWit8tCXr76sIAYPSzLzhQ4g1VRInMMu5owYd5vr7TjENQm+QYUXz2IrxEXeY1mYYjbLyTEJ0FSj3IAI4qrJd8u2Xc0Y5qO32Gj5Ss11D6o7LIoF9X0h1mdmYKqzd28mBg3N3cwIRIgjtFvNLy76JWDTGT8pTk8pp6ZgjTfD+X73MWMLGX7wMDL+AZhPk65XuwIRoAOzG3ATz76IYATCldxGizB6nTQRvAGrjitjtHqGFQ6IaHyiPWVjzV3XMpHL1sI+9cjzfaWcPbC+SXcFT+Tb7RE39NXuseo8KkGPky8OYRuPLy5ghF7DsLhMVn89pH8ubXbOrFCCK0HyNfOFBPQaIG8N1w2NbYDV9Jeusv5UMJWS9EdGr7g1ieKbhcSrNN2w7aCNDGCYBdb+kfeCFEulxtA0iul/hMiZk0aHA84/wATbSl2YpxV1do3RpHbXI+bKjEMH4s0CCjD+J3v/UhOh1PT5kTbq2nc1mMvgYqxTWWFBvY1GYEvzQZloLufLgYSHnkzIjFfyWsWWlz112jH4k7PI0gCgqJNNMYeHZhiKK+Zmog03u51m2kPWERLm9dB0ShJSlrKi1Gpd5woQQ45qSXpfn/prrCqyckwYGefQY4tqy4Xs/aNF/h9Z0g8XeqFPANkFKMMSa19z/EYlyvYYSBtDoytSy8g8uJfEGTv3IFbRNECVAQSx1JR/UrryOIluHa/aFAT2DsyyPKGa3XclQ8sWZeukIGidIeFsoi4lXcTqxB+1BqzKYE8/wAzLpIa+TKs9N5u6WB2dJpKl0HaOFCKSxm7A6wBqWrCEFFPN/TttH8CxTR6xgVR3JRKlkpOasPql35cB8mfOmmdGO6gy6WUztKuiBQNvo8KOsQnG75xB17S2KEo3uV/4Gge88qUHqxlNdGfmyya61rXdhrmAyvnD6ok/wB8B0gBuxUN+DR9ZvFy31owuuUAO+KmfOW75ETjLU78nEL/AFF2z5EHJTzxEKmxWXcZgQpYNBLUzT+bLwDHVZIgJyj0Ccsx4Gstx3ij6yCLdDDLG49IXYnAxaqWCWeaugsCGxjBUwijlKt6z/eN1QQ6U0PVjYIxCuyDrDgbw0j3V0XlhWLHMpaZ3/7hZSBPJLfqRFBpKuYcC+0oLioDeUoKLXHSUR1gji9JM5gUViPsJgRfumjmFet2rCvIOg7EN5mngQWxPvQTClLY6SiUhmg+WsqjAYAgi6ozENPARnQX3hYNFJUYwFALNdno/SdMmnx+kGinAcnSLEqA+qn7JTufJHPiK5BMzWgG03l7gJiK1YXlPBmlk8yXm1V/AwxRDA714ZuQSUWN5uzia2FkXTCOgvmYjoLbYGkqWS2Bv7rmNpXQXUhQ7WRZzQUpbTB2wY+lTMwcPp+oQI2PEMypfeMTRl5l1IqX30IoEyX7ypyuTTuA+/nLSA0Uh8NYweFaYXBIG8rLwIv54RJgo9SmFe2XIhMvOQYRLJqwSCxhW+W87O0tMoDWD6Qg9tfDmU2d6mRNOLh1/LmXC0rwg6Djq/1OCIECdqhswsI09CZJ/NkOkdgxNLICXcylDBSO37ZsgNzcD9FkZDvj28MQQDMG37Mq0PjCZ+mZ0D8seDJtjSOeVWLAWtr2xO+ASKzua+sOEHxAP9RHRLYItUcs83mUPOVn36QkGi3Ue6uPCmbp2azZDt9w0YOuvaY4M+bG0t1xoNUBo6s5EYTQ7ruawMDRRK7m5cg1r7TDFNifsgiU/wCSyGD5m8XUW1XPSCYcwe8tadoGAGi1PHHiOWhfSAB+bldc2Ysq/I0TTwABVoN48FvYSu35lUI1r6myYppbhHeaQLRf8nY5VqvSWSS3hH6nlO+kmniOKx1a6sGzGOT5uYmtLXOz0cYl81vXdK2jZ5Bcxv2HEjPKQF+VtD2jJLIo7NXIHd0Q6B/hBLPxm9oiCxM71nbyhdaqy3qesZxNHeGFLPlnZOkS47Ac+dt5wJsROSKiDggH1QgGAVLpJYsqY0iqp9Dv5y+vV1G/rKdGL8fHrFK4i+337QX5Zvc3i3KLbv0KCE3t7ws63Ips/AB7sDIWr1ro5ScAcv1+81yWrML6MLBz+CPeWDOiFeVOvDA2YA7YZcTEugdvlLV/LgfaDnFXVvKSwc6w7/pK08M3AG16m7ynZSe0PKvPFrGLsLGKxA3Y54tx/mixbFfRG0YErM8kNbGB0lr/AG79G8MkbrLbr6JeXH3a3lWYYfvQzKuXY3exE6D5BdoSM5ebzcyhrPA9JV5pFk+kAWRbwVadekG8sMp6fZB12dPnHfiAARHRvwqnssz58TzZvj7kDcZVMEdUntPtBYg0RR2lOVTTsPhvAd5n6N+5A1YJwYtEG7HewsHzt/KUjTyfTQhLBjCPeLsQ0ll1Jo3VWlX7+cFVXdq+3MPMxGteaExJo5QZjyXI7BE+St/H1doE6JS9v28J5kJksBI6H/YKUw19pxLaqdj+YDg3MI8oN9ZYGxKAL0zvnxFcs38ebeDDeliMJ/qrcyWIBBXnczkItkYDdi0hFi0c4fLi6kEWoHDp82BGA2aewRE4FKMSoUJqiydTFqpT6mlvK1IyFD6uYvMlXGzdWqFtYoNahcsd+LX9QStINcXo7zFk6hh6AetNDux5duifzEdbIvbtDNlm9Y70nTKNVwlEY2ETtT6I+GGXnTRkUGe6zHNle/RBa83rdo37svG1xb+kGULNkvfENHGwqE1N10Mdhi9WDZ0YIVdLgHioja/Q5O6Y8aR3H3JcVGg2vb/IF3lPUfaZ/TIs7nEKHpATIqECOqfqplQXRPhtGCgt0JKuPWy9mZhPn3BsdCeavG+cwcjPmDUAcOj/AIg1MFAbStRR6p3c0ZtsaHfnNphwZklibnXoddbdoR1SHHk792IY5BtKIxPh9ZvBNHyGs6FEDq0iJVynPf8AwheaF/WUvMos5P8AkHiAZE7nqO7KJURbVde9yjJy6NYh0g8w24y7EsYfNsIlxZzHKu0DL4QMLpuh+R2YCLNFZ5T5YIZ0yBRKCcXizVjswG6v6El62Sau9HTL3gi572SZZy+CL84JUbmYSuszIfffyhKcMiZmE6gDeHHRiS1aA/PpMvNJv37JkQJ1z12mKldsUXU38oIufBobYgmR9cuhCTzYd5jFeM/L7TUMyZhekRYrMJhAUBTunA3iTFUgt3yaxbxFGBwtYJ3wYB3giINA8AM0J6vJFAkLFbrrd0jovV3sJFBNQF+Xt5Qa7W27oHidKy/Qbpa09cr5G0BXgHXTruQQju6onJmPcrY0/mWEiUSNi5jfjcM0W/0ujDD1Ys++0r35u73YYyyWVLR3JVNzZXnmJTog/wBSgrcLQ6r7Tm09Z5IaHgZoo8bzMY78wOxaHgvgQpCYunv7uZYsocAfeGtO++uY2X6A1PwynWbk8k6hqDycSqUqMCB1wWM3MrRVKherD0DMqhdA+Uy7K+AaO8TU5r8VSoFbKsr3YB4wXI2yQ81YLh/EGOG0HtBWDqbyvbz1PSBdQuvNzAanQErGXCVlVhwkU5mO23ETkg1MDGZ5UzIBQNj7tpWCmKvzuYo2AKDFrPwqxBxcMvV3ZRrKTmKBPJjFSm7FGxTc94X94iE7PEOVA0wRn+IgP5jGit0eXHgURHR4GYmCmqmUNMOFiSqq0r7QLoMHB7RvGMf6JQ4OSl8EKRx4QBUys5EChr1Y8QDqGmhMNhw8u0FdsCNJ0R/xCAAYA2lMSiGKGJob1xK0KkFBviFaWgJrwDbZzLpArq0Q4xqmAGS0B9ZTiaaIJQPJ76wTmMXMpTuwYCyt95cRVqpLrljLUmBj/HPGE64BjQIFEU3YQcIAoixF1GR0CNlNBH2xFS7kbdqhm0Ny1xdNdZcGuR5x4ro+hFNukx0PV/ouJDZGq69SdDV9oS6Yxg9hmVE0SyHgJ7fhPAjtl5S2jcL88xxMyBEUaI16OrxdSiWEqNZpMW6DTcR75dhtnFUHEAg3kJbFFIfOX8FB4OIIkbHOIR8DiZqQe0TQNJLKA6lYTiO1QwuowVx3qqvzMN1/hdIDQRglXLYL1aYHSjjLvliUhomISU4bQe8t+7Lhsy9kP9CEgI6eAlkolGeWepicA0vR7S7s9S4PrKDUQRt7U+0E052QwcgXeNOk1j4VN0JaR5Dyx+YwBgwQDvEyk2T2BEAq1GR/iCjNvnLrp/AgOR8IkbNvcnlLFRTlFf4gyjrtuYjW+FStIdJVa4lec6EO3f7qA1RHVMh6kfklR9YxNORT6scteKMtKltr0KpTblyX5yqVTTpK5SGclqIeiZGXW/7Wx95ZCswfqqxLcnwlGHesIr35gGYNAlUqieYTbv1i/LG+7JCLVHADlYspxZaw4zLspJQADIGj/Zr35iuBKJ5Uq5tg17J2pA37gBY9e/WVKo14uaJcShc56+0rAFDFEpjiJCshtuDsKZdIJako4pG/WU1th1WO+ttUJe28tMHLKoPw2ekozKr1iuPqCtdkMMJQdKlZKulbaku6qmZUa1MCkl3f3hQkCpYOqbSopVomlQJomBDsCjZj4wLuggMrRHpctTl0y3zHqVt3BNJFcAe2JZFfQPYFXEJfgy4/YLudPC9vAKGcq4IthUIHETaaJF6TzrHlGQ7b6kj7aL8zru5hBDKlvsJnS1I9zH28Eh41lHL5RXXTO7wmaU8fnO+sHSWadATlRHqiXKfsb9Ssu7f+SwlQSnj8e6NpaytWMTN0fVGotDgJKhROzYe/SVpV30OI1679Ks48TG7KBon71uxRg0mmexwIjY3ZDoa9pjEV30PTrC+r0T5qCSFPEHwsmk+HQqNZ3gz4cphrYgho6Y3f5iKe+9iE27StnKjtjuOYeD4HEUv8UCSjNQLoS3Ftm0JfH+v7zMTAsOA77SxMEyswOqXtKlng6bRH1cHM7JbUvTEGVjQLmtZ0RBuCQ2PKK2cZ3kGtcQz1lsYYmcDK7CAB9EQK1vTHdnG95DE2Fp/EEqDlDx0850vSfmItH7ZUa2S3am5947hPUe3LNbeoTumXKyLx7wAqytPK6lvXWe+zwzXnhn8kp6yuGGdGP1R2sGyGBRgPHyuYUPXEvwJSvp6YmqINkP5jMPC4eB95Yn3b68iFJh1mTjpKBXBzMBKfn1lhLMv4BL95vFoeUolfVWw84MgN9aDhbKe4bPWII9fO5yQTRw+FbLiugsr/AJM8SpaeREdPWpfXOXrMRcqoCC7KBMIubmh4j5ln6AcMMpeKYL2S3X2hqQ2jpCxT5DqiLgw5g6c2IAC5z5SWc5lvgysLAEX2BvQpCLMm3ZfYxFlhlp+pLItR4XFvY2JTUHl6x1MQOkj3c6SjnzMA1xwdJWJJbhEyjyYoB3rUmm0i7ybtO/btNUTDGXhIpzWTuaTUStaw+oHmS0AM51+N0hh8OSj0hD6X9ZTLc3kB56QxQAWNHklqxv1n7o6QUD3TokZmDBqekXpwStwM9eAhzAtow+96aQsDaFG93Y+POKnoYmvKn6GogY3ZHI9VF9nvNKgDFmSsr1JdbF1S8azSajnY+atpb8zTyRtMRghgptogKDQynoTHJ6ouo8Vs208yBAPALuvzaawCxSyyfkX0isihAG7ELrw57c+81Z3K5TlZWW3R+jMD+SINAvrDSTGb1wcTZ6/vjrKYMhuk6wg4xvZhrM5AFJSPT34CAi0EDrI9h+YkaQTaAZQGuIWLcyN9Ywtnfno/Oa4NVPzUJZB3h6xeQbBquCYV2a/D0gkzKA2i+qspr0YQnrNPabguhWFOMyik6jzCAuzlHoNmMw3OJnxUPlwDnz1B47jfwSwRQURYYSqMJim2lw84NarT89KELed/rKawNGp3IsGgWuGdMxwZxDyv26da2me+0X0BBjpGKMkWHcFQgZgXAB9ZZYi9nmS1FOTFV44NYdoBk1Bz6Le9FiutvY4JWsQYK7SlwisOsURgRdtBnT+kHKLDgWnYNTNYmsaw7ZjO9xGjrAXlGb9rihFpzHRXIxoGXZa918MoA2ckcj6kxszzMrw7wN4kCOAvnc4yd7OQ0ENUMsHMofq5OCvRmvIaT/Aymex3jaRAOq9IuvER9eCahDmIlcZlBlgcLVOUgTf12vAYEm2fhPKMi2hP8zO5wDcoP7FQ7pWGXed+CNH58QcEKry0Z13SLcDXl1UdJ4GZEuCIfkhOnx8gMXQ5buO9o61X/Eodqxp+ImwkkaihhElhDZx0268y1mUJJ6ndnkhsGl9Fdu0NQgY622htWRcnBFL4U4HrwQZy+wMVN5tQv0CfO8MXavBQ1hh0qDiFyZkabS6BuSup2r9ZRlF7HePlwC2j2XV4JhlGtOtn3glwPopZVto36QLXg3apTDDB8QhvoG2O+8bTFGPyDB95jh93HUt5TuzMcVDfHpvHl9oxT2j6DYgol79whwwUsmsb2lm1VuCIhS7YVCxBj5P8+OzrmWTPiqRo45lTlxdHX6xg7pMfHvMMN5TKuVgomSnOHWcw7QODMfWIhDC0i+YVnT3ldXCL6GfdiFAOfafDOxJQYOo9rKHTrBoav4Pyg5hwB4Ndg2GKPEysB2QOXpROfpQ7izqzdOZvS/6cngwwYOmUcJySsIBz1MDQbL3OWCaKjNERXbWg8ya7zbuMWmw6/gIGVpK2e3pGW3t693SYofzAXiGA7b2BKUZZsOHUUkqnFvKEQKbnC41xuwCdY5e1tsOxyQFx6T8GO17imjdXX8EojIMEDjKlFnd0/aAQhqizUzNcs3OW4+9xAfAjTmOwdx1jWwZXKurKfCwwy8GxscjcASXqpb1dmLTDtcUXmdzKam1pdMlHQlB4zaLHrUHhinmqDzy0CKBcbLBdiPpUFrHlV6sLeAUnRKuHDGkIzsiUg0OHQ6RJw0ohSnpbpFf5vy+f2heqBXA9IeCpKg5g+QUjH4G5xDh6TWQMe1IIxmquHlE1gUZWyumr+XJpl6OjwCKrWaOSBvUzB9lWIGfhzBFU1Qb5/GJetObyriAgFJK596Alao1lB2HhkViaL1jg0ZIRAWx16XxHNSKboqRY8uZ1VXeMt/VAzda4PSFWFQG0rhAlCM28IjKwFgEsEXC7B0JiFWlNSrynZ6Uy6ehHL5NWtfzDB5QYhiALvjrNWpKXVuJWirqb7jDTFKRmZI1YqJVXV1wm28BeUIH4oATp7ntCXETsFbmunMxWgG3LzKAgYa2ZlUeBH32U+7pAkO/9UxLZaXl+swmDNl28FhbF2VF7hOiRjCW/YzhsAaBKxDMmGpo1vG4Q5YzruSWBAvQhFJRVeGsqyIZHT7JT8uXC6MMVE8LDXCWdwisEuSjiJIhNq2cR3bH06Qk49HlB+1K1f7MxxAiRIVIlnEuYvVL/AIjtkG2kXeFZ+MQTgtyF8fOYHY0Q1dekEIltGJa1PM0KA1dD4GBbLpZp1lgNCK+TAbPUYaEG7I/3y/WNmWNDTHPdDHBYl3PVEjLGSI3siX58zSFIIogWhhtcR7HqcQEDo3+CQA88Q4Z8DDSKlWksm7wx9wmytD9SDoh7R+kDLBySgo6UqQPJMtcRlpEl+CJ9xTRS/WXmO7yvPwCkJqtY8mYcXNB7DBFfQz56RVCJ2Fur2lVp5PvMwBEAhFEIs7SrWauFFSmrM/SNogXGtqK3tdZWVp1Y8qmm+JSDWKrsv8sLSiHKLRzOF8pXGBaukeY63HoJ2FEuxveP3t5a0NcE8Y/jlpCvkb8jxSpV0ZTlx1lVmxXslEXnFtEQsl7qcsdM20hn5ucVfVg5lKAyuXPhhGLznxzB7wtcs/6E4iPTJiJoYUOWX5TZRh1epFAp0irdKMABwTBCLGZXvqG19ob2UAcmZp/gQ33ZodN+LlwioSTj3UDJnMAyIEELRq+hDjUX6vj7RijRMeGmWC6kdeI6RDtH1iKGNuj1iodMYM2H04/3LrMmtsPfEFRz4C0U0EAGKMxdklCNJWBSI/4IjGg7o1+dJcTfb0rEOwe97hCYxSnems0iRIIg3gFo7kQf7J/tMshbpVxzQxV346KloKZq7uI1pQ6klemfBPBBUakd4j0UbnhiYe6RO0EMRE3+sRXulzW2zMyCa+cqEFCaVANTELZVsMcxbJcZC6Okj+oUXv8AxDPIvrJZ59pPaaO5hA9HmVS9URzGzqENRixg8/Bt0jaUQFJKQaxrcV9ATQc0pqhqG53feZJAaHD0YYodEfQZgs9ZUhyEq5TGRSaldAnduM+zDcF1EB7srpXMcCi6m0KCVaDVaC2GKg+buheE4xB0jl4DUklV39YivwnWVpBwCWzLjmPaAHO8wcDz0iGlqC1CRhOERzTKF2uvSzNoVTV0eIFmMDYevMMlhkfTEvPAHFFBFTqPSYiGn6OkshGOuY4MZnFhjpKIJOqAbs4iqeVq4dgI9tS9eLF/2ptkQmGgtoteTp4JFVFRHZyQ1ADGXX8y4aOuldSxI2yPUMXx0DOnEEAYGMo7KPA4DCZDd7+BVeHLkONy8TcPANXYm9Gv12gKoD0b1nBn6g8pUm9yJzNNBi3AN4dWacQ6Jwkg8DxwzAsMOlv+TWQ8pUDkXJqeTNMN2Eq0fiHS3mA2gAM6iOUqsB8kyrlRLao06wsspiF069JVK8JkU6gqaax1XdhSivVGIXdPJs+kwQaB6BdGzrLwkUo7qWAFkGR1uIDDVqEekufRRhtf+H+rtG6PJxTS6++/59Z0eFNRcR8Or0A18QGgv1Q/EZwAHMCeRldGiMB5xHxdrwKQF7I5N7D2o94DQgbd4K8WhsxOav2PzDS/ExpA4OrpH5ywt3R9IQK0LZK8T6UdUTYb6fOYet0eh4YYFiGiQK2wHyJ7eCSotxKCxqQ1fjmety10esIlc4OMFPtvSUFcGyTgj7YW90PSGC3b7Sm7iAKNIW0IDBEuL6sSmw/MqoajPzR279IrhW3RvI6R2iR6S8gNG3TcZlTFt+8eQUcwrvG3SPgcgOWDD2geg9OvWBG7qXe4h/Io6QIp1yw66ypVbWzdJTTfJx+DKed3QS4+AwJ8Nqzc70M9X4TvW7IYioelv1JqJN9KfSV0WORyBHCW519Q5g8xvs+Zt4c+U7zKPKVd8DdiU/EZgwOh2dvxU1oQfuJe0Tcr7EI0C2LTpcGMNyTcx4dk1XJMr5hNOjqlxZCHnpOdD9A+QlKoPIv8RD0VcfQ0IoQ3la82X/oKaxELo+qbLmscTGL1nnqcuiCqe9AyqI4MZl7jDFL0bVvE+lcVp/qYIepfuN4gufiofQT9MiBb6oA7wvntJlnwcoHkh1oc+g55EIqMZJkw10g15Ma68sN7kRrnViCw3dvDpNeHuQE6XqJwPWSsQTV18QmQLBhIWRSkz0GDzPkSYdZ1PWDNnDi/xj4mxz9yXkUb+tYponQ0HgNkQ16Wq2DuezjYlgAdTQ+GY+CRu7LqI6ClcwFPLt6wohYKneXQdT06TDxokdoE2E5nzc0eXpMmWGATy4iy+aiYVyOzLbuDROl4+qZFMCtFQULd5ekLlzLl2G8y5sn2ZPvNQ/Fmn3JoLu5tc31iNU+edCC03SPKYOdqF8o2oDh0hpCq1eRj6RtL0+vmaKWqOeJSQFoXvjJNXUInk+ye0DsFrtIpCW+qBlUEEPDcj625tzgHbtiVzmkRpvhCz6e6g0tFWSmXT8kqEGwcaMMVrA2dzwPT3Dd5ekY61vtuhLGVA8QZr3JoVPCMXmI3Hpp4lBBG6IfvzeUpWGwaMOsZpRqsYwtYj9p1hiQ0Qr0NDy5gJW+lHhRPCMZpyVWYglp4PJ1l0athCuHpAJzN4dYOTEaWPID8w2OWdUcvgrbhaNvWb+UtDDo1uQYAqtY71KQIKPcKGkPHc7QvUveY3biY4hjDylIqU7UeIpRJpLj5OqkP8IkuDTRGJsTMdkm6kqFPcRks0m5QE+7zhwaaJFVpUGwbVikH2shoKVtKJKpZKqfkb2WROPGj9TUzxVniyp4LyceEyJReoii0BN3wBEVjPWOYZRyiG7QqdMTMIcHvGMnLSqAGINiGEafQMyXgdXyFyzXh3IxCHmbVt2/rHy8o1akvebieeNA+0d/urUO7Gbnw12QJXEGsXGsup7fHSDfgs1VFTS6sitUcHziVL1clebYl4USr/ZLdFZTHUzVMx1rCMMdJl61jKAuHY+GIOjENnY4+8U5Lcuv2jXFbBrBRjq8oSiRM0za2I5gv0KIQrEmEYUwlnU9kD3NZuRKnit1XLLC7c5MrOzn0PLBrgu88S/gi3mprGIi2roEIAUMAeCji8bD6Ebfi65fclsqwi7bxaBcm0Wsm0970lS0k3naO0xC89qkDqQNL5hDtHoyPBG/hICVS1xoEzgoyfAwHwU+a3CGVuu6e3SD2bP2g6yroTnQTYbmEYDPR1jeE2+2VWpw23GkKjgI6X/YRawSbPUdZdgqvptUFM3310PtLoAHoGCX9L1hMI1E9kmOkpgR3aAlpFCzecRAmMkadAFY6TKMeU5CGSUF7cSODZNas7kM7BMRjj5duBMIJfFxW5uRaRXFZSnCUTwAQnEVCgUnpBWk3DfYirQNRpTCsA5YWBSyMMAemo8QNVRomVG57XV4ilisi7xjjYo28nWBXqhWtw9JX1YR7WKH8zrJE1XLCkfAWU94RYN97GVAU4mjT9LR9Lh1JqGxzKpYt/wAwr3QwTsHUrHD+xHBKDxUlYZdMQ7S4++V3laLR1gMuwGewEoTV+Wt6MseBdfiAgttd+rAAFHgeEqWTqthsecpK3ABejrNa5GifzP0kE0wfZtrEdH2zzKjMIvgQ4vUiV6Zj5xkrTttAJKb7sMvAGJpmGCBBoxVq1uyHKZSTzsDeKLWBqJzbidJPP8Ih4aR5TFUarfchGPgZEFyi9IL9UHWaTPix/p0jT1tXV7y6Zm8eh0ikOlaQT9pLkA6EHLCTqyi1fBqvAaY1mVL71TyRwgDbDyxxWysDQZY+t1Ftnzj2hJ/O/mA31gJp+xtbp4ggSsRiJY6kbnPs3b0mFtahRxKt1VPRpDqiClat2isKtWuXhvGUC13ulTGg7P4Avr6w79HpMLqfcv6QZYVHR0uGFFVMwgql87QWSq8wZyZjMVlDtLQtLgPRf3pbd/TwH6oAAO0pkG6N0iHGlZhuCUQhBAI1YTkA+tL7XjaSoZHmjKej5RswDnFM0QWjQIXS6u8GkQphVEC+Rqlj4ttQQ9JFMK1Rho/eM4W5roZV1xCI2DrgSSXWWNneUu4x16xIjm1aj8wXV+J6CdWYRPAslm1+AwO5CqfAF5kozk49OJWKDiT6BTVKYGrtTl/mBwMwEDGIyoOJyoRb9IVPVJNI2Gw/TdippAekHCWOMKoYKaZ7V3eCMxKlQT3/AMidZmNXeBG48Hm4BMBzuIVRioaeyJYwdi4lbOIAeFeBgggsmqT2odo4zYVhMQGprUH8tXNG0+q0g0H3n5gQp6SvSMOcrPhYQQpm5j9ojKdmH1xQrPZYZbsdeIlJXWIZPtlMV2JUCBCCNNYKIA1uIEoelBtNKMTC/XwdQA7Ce0A1qhT3YxC5gaBA8BKlhrLBwhEZHEwiF0bry5hJU+yjFgRajSX/AOmUAe5QI8G6m08AKlTtKuuGL0Bth1sC7QhsgpDN146SwNbAbHBGGe0X5gv5X5i/5X5gUzUL0gQIEek9LGXcBtwjX0SbBMKpJXWPSoQzruYcCSBUtoZcZsFR6G8K6iAceEajseNop0DKkOkIccr0Jrs2OpPAqktGtkP8JBfmRIGAmRQpZGaI/SOmvBvA/wBgnRYgt7zziehiNWHkEjE1keJQzRCasaia2qt4HaXdGxFKpRzfnETR/WsqaqjLLFNDZyxJZbzbYwdoMPunQCCbolxMywoNa2XTEC4reF6XPdFamrGledv3JjClfcQ4Bq8ziZQ5SfpMXOonhJ0x7KMA0pkSpCDCCb4o7r5ME0B4cnJLNSyfabSw5HE748EiRKbmjLZo08TSnBGKetKMPfqI4T8Ql6bVD3amcFazqvxKBDsE1EGElQXApYjuS1Ze02f8zcD1pAXv6RVkadL6kas3rxBnTV1JgZVHJNYxXgabRJV7QiRDcH9eJTL1YXEYmbhsGUrnz07yrY9lmPEnSOkGKQgMrYMsuqPVKZrSe5GYM6AVKIFwgjSa6RZbpGs6HJNICtgyqExjTJJpKyqGHsaUgPs/T0YILw1KqWO8aqOOYRdyyIg0Yt4omuqE9yOkfUswFuhKkAy2Alz1NdZcvgCBHGk13plNRreEAIPDS/MM655awIlejB5Spu9p/kQh1g8VUPSAQKGAPADweuJkBuY3eIICdQ/SYlJ5T2h5W9wrMfuYSavnAYHY07ml66fkMJZTCG/nZUVFbNf8w99fJNCAqZIakS50s7DyRx6Qa7ufxLwMUOhpKjzpZvfn6QHmBEMYb6XVMEeXs1HDpNPbx3lTJkOWUYUD1xGQXdboekAER6xwB01TXxGjMO0dm4uAmpR2EvfVwmj4zD1lt2oiIBbM26mCjc9tVmBy/dpXAXBp0sMd8/Ulo66IJgb8runSFmKYFxWioGQJHmGxDc3jgvNbuUuG1fWOusoQ6Oorns8wQ53rZjD4BxqyjrzGAaEBmD/FMNZ2QUHz7xfJCK3ZUazfh9II2BYmjO/hUSVTK2Qv3iKw+QQuzK7AYb20u+8M1fIY8suUaacKhUS2Ksno8GHwANiWTHpuJ7kLkBajF+GRc51p3BATWZZC+P4g3IxprhLIlyvAcolImESIU3O3yhtBbBjFC6SUqdnaZXqLeQup2lf6b8kQ2uJYEJ08Gsyu0YayBeK25meoGRk8QirmkULDT2CaCNi4zxGuq/wjQFdlm22Aqub4NNpMKXSiYdaEU5HlDmIaeY6fAPAQldWiNK/6QckOHuvX/I5nYqBHzJyvrcZuqFTEIyHZ/MFMMy9zvfWFJZ4GK3hvR3iXzUt489Id3rno2+cQVZrYLCU3whFxLpBchUS3YXXC0DECd4GoK1bSxqu65YzhwG1qWa1T1mue0BmM5iuZ+jn4cSpRXuEOpByawApOzfUPg7CEuwG8UOxSN/4hqllQ0IfGjdCZMH3UGEFwFukvt1UR7r9pQt/mgKOLBLXr6R1ENqEpOUBkPoqH8sAim6uiPzNEDve6OgGsm9UKELVeY1MopHeW8r5yERRqnIukThLUpmXl+Q/zBgWmq3dl331PzBxoX1TRJJK9OZxwDW8Kp4VZ3lfppznBJ36dpgeozs6iAbLY2mCbvTx3cwiqFgsRXtdgSLuRUkvf5xqWzbIc5Uww1sJ+JQIRdWlYnJA9ttHd61/e/MxL8TOYwL68IxWaLgNB67zWkQbDGqVdkGYqfxo0KrEEq5tHeQuxBBJZlAvAAUVuswZUqJKcGA+o4PdJo5HmbDzXw0ToQQ4BjPMjXvHWb1ubcr1fmdYS9Gyp7Jr4MYYhZofrxTLmLAkfBbJACMyOs1sfUTHpc5Rl2icU16MHobb1+IgXCgGzu4YRglbyr8BdAFq7Sxuyqq6jpNRr9A/Mt2hjNEhYcb4WbPUwQg6n/Yy/bp36PWCdnvnkZpz3YBEHwN489pjAJiongQESiUOrF/C4pY2xfPaYHj2tN0LPu1pUUXrmgA842I0aqwGdNgzgiThOaCVt3HaHbm6Z5OjKYQoK0jAxarGaNDr/AJmblXRTDLpPVYKJhVBz9eh/jINN6NNECbMg1gRd2s30MYKWsiQJjtE6skBy6ZfkrQNVwhC7GuAbeseFJpg7SzaCfkyGAtdAnKXqeRB9VUPzslQ++Z0YQwVwnKxgKfgSiYKWBRlaivBe/p2Ra4t+nQn6CfpZsDDSBVMQWm+3L55BokQq9gux6MGudJcLFDu4dJhIdLaK6DMHkzB1hV/AhuwUGfk7TVJGhhdAEsAz0nWwVWsLw1yFQjVCBuYRik1LtyV/nHVcsOUKU1QVxmeuvrHDUMqxGWWk3RyGWF7EOCqbSPZ003Rlwe66xRTOEl31IiUEoXNS5m53WdIcMPV8Uo59rzlpNVL6w646QUjkahSt/JLC2JlFH1OJbUzWNfSWUbRYg6LRyTPiIJyqV94QZ/SHp5OkWPU3Bn6S8gw9ItJXONeaRAm2Rcz1H2to7StYVLcRu1Ala4vPiM+Ex/YRb1aIGaw2anEwi8oVTYTRnnCu+Z1cS7MSpngsLXaJzKDx2EYgFSO8v4XRufEt/Iz9llH+kV/coZf1h+3FWx1gm1HkdTpNYK3mjrB2eAMprVlomj80WDUrx+fEK9GoxCX5YZsezgy1iW7ARdjMo2/yFL06f4ojZzav5EBAbRJl0jWAy4I2SL9hwQhqAlHEt82w90XkrwnDMaLhDjtFtle61IzrchN3+zDjIaK/sir5vDkitY/q8/BjdAKPdmbWW+12jJULshCMwcx610NXvETU5f4Lc16nQmcgGd1GLzk91TO+NBPxGgrUCBL+Luy8IpmARXYd1TG86NrvD4bI2OSNHAtDvywXQli/rBZULDlEJAVtD2ivb3T5rm7E0B2JRztdZUOQSwy9HK2zn1JlpFFTjw0QRI7fTvKTKe3YlxVtwTmfLYc/6z4jPkseKOpXmWY2l1GMQcZ3cfvBwAsSPWV6reiaLJVthvLf3UJjq9otsaLaHE5V5yr8k/ZRroO5KHZqIiQmSaF2lzkb9YmjSWtdwgWBtVKtcyjlLL0Yv+c/EQblAF1jf2hT90ln5iXJIuSPWCHpLXYqVwb7XAGftEd6lSxRTzI9LvNOv3JajFUK7TL8Y0Q/WOdkcQcgqCdy76YKEFrC/eANbk+iDIA6QeQkhF8iaBOkdpSBto9ocsRR6zSp3qyD8kvhe6etNSnd5Yh20Vf3g+aIREqQcoGMzxJQGm6Zzt7w5SFL42TCGF0G4gZnfyuFEsBeCnmzCCM31nRVXdCvsoOjLbuTT3j+p7T9TP8ACT/Ew8x3SZPxdH4lvad+ynAoR0eJlpggFy2NpYTgbI59WUIkB2WkYyebHR08I5L0gRZG4R9qAApGpQyHAmMx6n19osrkCSztRFKUEzM9OP2ggCggVBAk1MDU6kNNi0sTLETXUcrl3P5MqcuRaDpLqfDRhbNrUdH8SymTXcRkM3xnrwXdNXdZgSrmnaA6NTC3nLhEBZ69/aAOON27ymtfK4gXqhMPBLvm5ZVsdRa+n2l3j8ZXpeDvEq62dPSLFiFZvQjMdK6VU4jlsRQHEsSHgubtSuf4Q65bEwxGawkiBKuuOPWA8FQiTpO9mm0caHaZ+w1qaDEvYE2XMVTGzn0I/qSsvP28gQIQh8AqV5XFoxlTPnpHeCU4ZgqOrmvMWMzxevdlLOLVlCEdASiB/kT4RFePoSzEbYekLqgoCEWEI0UUHSoKO6vfIgb263ZEvnoEIXszgE4gfpDwZseK7YjeomTcQgD0ECvQ0Ty0pglf10/c+6AKHYI8cRjSOBpLzJ7wy8dVMpUPfP38LM+pPq0PxOa3VEO3rNLQyMEeoML15nXoPgCEl2nszzwkx5idhVy+glFaIX3gnbrRu8BpU4/RK/oUV8p2/wBQ1ShgryxLTTMCY5tD73DdDpOuMSm0qRl+9pfiGu3Xdl4lvasb6gHfFcHEpjhxFBpQ1l/qX0vsNStBsWrIVsPrcr/0jGouDYFd9RxrCIiI5+PeY2tJ24uYHaOoprsl52cSklw3B38IMNC6bwlqHTmU7yd2LHRY6ylslTQoCi5r0SGB5qMgUXcNEpe8faBCpXFRJUbwQGzdpuuSkwln+M4P6QVf05muwOBxW83khz0gzmw+s6ThNbgWiP213ZRrlBKfAyyanRAjVt3a98dl+ctY9Mp5kq5B66beAQuSIDo3hLsFL5jaxRbsuCE1U1jFCmbpstIdMGrZG7TciRBLvm0ZCTvl3wcxATkYsrLDlLI/IgqxajhF6GQtZNZomAgj6BGYChbgQFkwmUaRYQUDGlSsPRt3DsxiVveZ5zjmtsOnpMMTt+UTb8TrK+M+sdeUAvoQKJKBCKlYjeKtbYg7s7K3OIqYDbSuXtOdI+RjwiXFeGwcqA29Kd6WrH0wswC2sTdqFFWwzDw64yxrzJzhnu8TANSM1Ne1juaRNr4ZC/8AjD/VJd/lGMnzhQ55U2IrPAovRt7xEEZLUvaRfTO+TBHSWl68SrTEbkWJdjSWF1+cuYWJc7ofbRTzvxKQdxmaE5vPh0j6imCBVCm0BsJs2RTeaQ0kSiaZkSZPRC+oCZVDiKGoOwxMfGEAX2AgrtIWncnq8AXQz5skdawC9I7VZrbJQTWVGL79pdGYMq4pMjY6UoZ/ioX6BGagnVClPRCCM/ZVeKB1mCuiNC8wLJRKojrMlkQTUycMrgOkjmaLceFVDHZHpeCJGBObM8kvfyL0mfmWePNCmjAmenSaxJXgWpt1iggDk6nPi8u8pyM1HJ5MoOw1TqOHqIwvVFAT9MMYkErwDcBWEZyjC35IEr3Y1g+ylhFA5ioCDjeZZjpEN5G5K4/1DvBSEYK/gZRixm77naI6HrdfdNFG1yXEkmpOrLUbGdM7xiuJpwdoal1ioxKde0UczWUb7Ao3KTZM40QeVGhlh4DWCaJUVMTGRrw/2M0a4mzutWFxGS5GSpRpWbPR2gLHxOku+B7R4K52HoLgMh2IGIECVFLYl648dJiZxUxLM3VOCIjYJUS9m0IvyH8kK/w/KPwflA9CcAf6mp217fEcukIINnXYjRe1mIsiDVjiLMRehEEy41Zel92DDGS7Yf5ufr0IWv62Sl0wN0IbNQvLMDgXGe1VxPSIEnO5SxXbUMIuF1sO8o5ZVXHluQ5cEt6/N2iP8z8R79c/iZsXB+CWK0ar+bQ1Xen4Y9wFTRxx43czTAvtxGeDgdbhtUOhCvdiaYqAej5Qj6Ll2z2/JGdVN02LPf8AmX3vv8xD8T+YhTWssfmMeFplS8zWU3TjaY0jVunxhIgOkMy5NBXtvBy+WaJtvFoe9wmeu8q6fWbV93+Z8r/MX/R/MvjCDD7Mds6GCTM567nNhWNJXeLCYQTw4mUG+0yRm32YbIHWBfnpGnUSh1uFse84TWGddZ3hiW12cR5iHkpSOTNGvWbUMt7pVChOkMV4HnwJKguIKLtDSUI3pwfiV+j8JYX8naHU7UVomABfOYSLCs9d4ZgigYxWakLp3OPCoxUYYaozOidvWV9rURLBneaCWqiVEhQFUAFXsylsa5RUfx7TK9ybnhUqaTD4A1Fkpy1/ixC6LZl+kV0wx+eEAWqjKsrM3tSK9NM67NJlxaOE7YaJ+0GSGgeJUCmUZxhskBuwaX5NWK4W+kfvWtI+kmwkCMZ19UBWBFO/qYxdPLDsIaElBtCBA8LN0BcyzB9ThOjqDtRheRtp4j9H4vt7zaXxjAFWOKlXPbDOV+bwUG0zBlYNiEVFCuAQDMWBMtX2B6TVXrWA7TnDoRYkjo554rU7hYNkFyYOrI2X2EpBQWHzf6TZDQssoZTeub2i/qWZpR596R8lbpj0jaY4IxWUPIaylqdmskNwpzTW0DI2vZnvk1OV1wxHoPQRCiEa8UAwl7Oses6vAygXnp3CeukHRCcL0oxCGhWJ75dTSY3MLzQVaaTTM6sqlepG1Qx9ZEoKurC1amtok/RgID9ebl29QWinRVSomge8alFrIN5lJa6MWHpMNyCBySTowkoRu0w+Cxjr7s0Yx8IpwYJczG+Opb7S5wr5e8rBeUhhLQW2ZYwsKeswb3hG08gUSiWbCmUJ3GgY0LkLlGLdwNiMUIKG5l7cEsabjHTjG50RPFe0DQ2bPaO35pZfaeZAh6Q5QGph9JtEjGEPDB6WCgdSOiDG+0I+q3WFnBxwmn+hde8GgbgsSBRohajyMS6RLPrAV3FofOEbBOkYYYSUaS9rdaO+Mo/JKNbJS2SrBF/cBQWCXmQcN4RTTf8AMLr7ztKXwJcsTXxVqNbDHYZ8oiUBn7+a/ES/OPFEacPMv2hChxFGavMY34EA8QlQbFXeBIT20es0g9l3g0sV3iqrgxEZh0H0lhg8IhY4/Mhm5O5N+jN/QQipKAgSoEU+m4aDvNAvM/WZIXdZmXocR+FT9UMYADWogJ0FU422HvKPyTSA7xWkQXRhMhKzzoIawwZi8tgMG83+JfA9+ZT5BvCLNttbEqWz779IYDauGD5UjOAlCFOkDIXaGdIQDR32h8Et9ZvfwtG5dbYMPvD8B13g11cFdQpTzFO1Czqg20D3r1mBFc/ZX+xGwjHSTTpMmQpEJUFpiaPDzPzKvHJpFbQEAHSHCNoglu9lA2aKezSGGwN0GMkNSxvHS66RJ7HOaJXEBd+U1rNwlySgLh/OW7OKvJDTOsHsnKO3zeAj2brrmBT3J0ytwzIMHstzWHEtBbS37RJItlKa+fSFJ1lBfq0TZ6kGyFglad7WGcwLOk3gJjYhvBYGEOHzmGusLRHEy3+GXWqZcMsKMg0iDK7s53rmX6s5YQ1nVLGFPSULtY1VM0Dc3HeFdMsYtiemJJih576pd1Rm92giQcQVirov5jMATGYcrlwA0Hi2A4Bi2BFQYuW0FvqvISj6ezEoEYLEpmG8AngSWzD0Gnkg1baAwOSbL055JZim96hM8nY0kvbQ0jiYVVVzJ1lAGx3IlQL8ZnCVCaop8+eUGg9oh6Mf5OaBr/E0TPCz4BawSvEvMeqqI5gdUR2pbowFAF5SVZ3gEnlF4HVZ5NyGbq9yJ2vKOwr2/wBgAi3hXYQwo6BtBXgCXPV6EWvalDwapiORAC8sR8WqvytM7wuug6Ivou6JC21d5d2Y+iQmBHrMKVNaXaYIQItToQxotq7x4Q3O5llOmLeUOnF1G49TJHMZB/3pZxX3mzHnFpW8/wDJnLubeX59o23SOP8AYaeg9EbezHgNaMSLqLgq8BCALzvmkSXScOG8cYea2RM1LdZu19Yc67sLrPNmORSZfv3hfmCQf8f5Sx0Gark8RfqViQJq4Y9C8MbwMhaDDsMtpVGCaQA5SwWd009C5jUhCx5kWrTcMiIVeSHaPvnFYlzL1Ea+JB1SlEGDRZ3Y8VBYxPPy41pojR7gLg6UVJ0mjBosacmWrjkLLtElxYP4h5XtdIFyVLS0buhoElnfANzG7CCqviB7J+il7ygR01qMvByRsy+eqeU2gH00e03Bz8zQtGuwbdopi50rMcTXfhm29kem8oezDpBz9AWOtQ9jOG7pKTomlqrjiatKIkWr6npCiRwxPC0NCNiVeqjqMI2hmL+U+YiuHlBXk2XSnbOJxEFqI9QIclzXSYxn1CUCg4vqdYZZ+Uq2MMfAu1RigS+6B6iFch5y7W7w4Wdlo/WXgu+QFSK7x8lmHoIFmoHIzBpDa0tSjV38IwhZkiTVKlZRPVfGm2Ii4aBZYFGXofVjjcx5bKqNpUqVAQ5TDFdsb/gRf7W1nZh3RxvD26S/SbfFNam0F7sE/YIb0QIFr1gOnFo+5EfNy3Z3kLIGPA21NjmLEywhZtDWAnBJ6m7mnQgJJari+3MreihZELA80A3vBF8EgNpSaWQd+8tKa35zygxEhKGWKp2Ok6pu6TMRKBGmQxNZssxVsfKLyJbr8YYW4iPGDeXKILjcD7BtGS4oVKunVjKMZX1kEqNOMJdkguIlRGxBajkM3/eKDsQc9YxSZi2ojd6QmlvKV+cBTFPjabTlQafMTAk7xuB7yCr3bbafuKBnNd4yIbK8jMCDp6QQBClw5jhvSzHeoNzLSCDw4lNsFMY8oYPZPzOSPjmWypGrS4Pei7PWJLI7PzLFV7JFVvqCkyDOE5v5cuxupiRkcdDQg9MgTb4rOsviKiJl3nDB7sGkxoy5ONDew1UG7gDYt6PxMmph+eIPR9Uo/JKeGRSGp0Fdm0BrbubmzPNOdGXyeZeglVrHE0VQXHEJP5M4fKLFWoNzZhK6n0lD4GGYxC6s7wegAOjyx7i2uF1g7XGo3JULWZaSmn7/ALRLlRumIu23zQCW7PUY5Mj2dJ0+O/PcRty52qEn6Q0MCm1E+XsljIWLQ0gx1P1MKq9LzEiSseAz7yJAEpUQn2R9HtGLx1Egi0O0Es3bI+sEBOgHcjgdXozYYaxtfdwBzDtOE0zqTu+dz2Q0FPaMbeAt6scGWVmWVNn0lkLakwPNhWMOnLc8B4ENPgaw64EaHflnFqfPbzTdhXXQNhDQOgwBMgBqvpBB0jqif2kB3fJB1CfHSa4MEX3QUraW7Wq2oymVjmj+YGI+ntb2OJTTrOm1Rq9CKuApvIi8ubn1JRVjW7O0wg9ITngQJVLcSM2DeAKig2iKlQ92bYa1Wq4mcsQHKCNaMTthxKyJvNjAb6RxNXhSwh/sEP8AJeFhvzkoLXk/MGW9T4OYjuha0JazPpBBM13c9JiEWOBitoI9FlTiaN5gywNv1jXRJTYyYAHVg6IBUHWf6qXfqJsA5yxlgoErpUtL+EEax2/yDfg/yFBoul1lM6etbm5No1k4ZirW3mCaCvJxGeyTMAzQImaJbzwSuloqeMRyemTYn5RmMVUhODtNedCmhKuYC18sl1aSpBrfKa/dkPMI2v3iGqrHoOkvoJV1Tg0nG/Q5Y+817KsV2nbrGgwar4x6QHy1gIbuuC8Q1v8AnvC+1Sk0lJOQrFmoxCRHJl59GOPwm2GEQrusRZ3Rplja2UOWJ1L2WVELvWO97yldUOhlSUveftJ+6j/uT9tLe95INJtT4Mocs884mzaCjEGEzB75dZbP1gxh74TOIYy5sFXxA3k5uJz/AA84O6eBgmBuqNzaatKmz8PUvpGynJeH9Iw4pYvWUJOnDoyuYNrz4EjVRdcuhNQqty7SomSKURnD5vDqsB6N5woUeSWlS5T5MYfNuQKvDa56S6Nv5QzNucUJO6tnvASdxr2lYlSjGzVu2lRUy9KuMm0PH4GO4EqHa+9lxJp0dobjWa+9nnzKlca8nmOT2yqBKWkGh/qW73f9h/of7BgF3f8A2COteii9G0qppIDeNhpTZwKeldyxsHQjoQhSgMj5rGVsuOCYVta8G7N30eZ8plt7QbTw/wCj/O0+C/Ezg/M5r0gCUCDmZqy+qNc7SbT3fLNx03SAcBg8p7HLzrR26MOt03uYubT84gvw+3hTCIAGwEw1YpNRoWccg2HdmCWpNRaoDaZQSyA0wGWdcN+Ih2RJeuZes9EERSKh7zliPIinWfO8R8J6yjVrC/JrMGWlZBYdh/qBLt+eZp+TfPWAoy4NJfGIczlWQyX64mcEMvmnM90wLEdn1YuAO3J4YiHsGO/GmKfTx1u2hYaOQpBWI/5CCtp2RLDeSMzOqjWEMpHq3+8Zjki9sEsm5i6Qq4R8gN8GKUIITCrmkwzprG9gipOjWUapDfLhrtQ/6cf9mbH1p+6lU2iO5uTIqwWvLSWbIyt9402qJrOJrDXzMIqgxAAsGE3NSWYU+8bfaLQS+yyv2MOn1M7H1Y8B9WXwfVjeLfazDW6MAyk+o5mpLZbTpEEWRVmMPMxBNgkB3jQQzULdxRKJteqPL9MBvhLcwQwa0jmjCcWyjmY0IAjq8x0Zd7cwEXjncmEudoKkG1mov02nJMeBiV4HSujkmg0wB2ZGoK+dZJ3ln8mu8lX6YV2YttdssOAopqYsmnLzn7GWP87jQ6zDGI54mo7MtCABfDRhcHfthoTZzevdBR0lrwlY61rxvFDdHI9I8xZsP8mpfDymaqfnaDgZeP1KvEyUxO2NIN4FjpGSmOrAY2VS59eSwguq3mOVdV4JbcjSH6sVGzSOk7Btrx44xTwABvn94FTOL/MJdJzVlS+XHmtkcbid3MPDGxrCXZNhZsrisUKFUoG74DZKII10L9Z+xn7CfsYL+WBCu+stfbqdM/Osbs1RYtjWSBe1NWV4W8wYeGL31myWNBletYUOAI/IInNOkGKLFehLuhLGFX2s/SYrieSPq/SRgKo0ANftM+k6VJu16Yg+o5VsucOEIPHYTO4hPrM9IbwEyTZT1iyMtaOzyhuirlP4EVL2Xuze+6NcHrDz0DDqmzFGpjynrBC1veLuT1YNhY3vC8soYYzDuJYPEevR9/aTWFYeWOOqX9fGCB1GixziBmXPDOk9anz+dYv8TNt9c+cmw9kf15p1beoR2wrN44i91o5IlYo2XL+aqZzznWGq8DaFME769/NNQsyUXgz0EdLDwI6WA9IbJigRNIHRKCy0HPSWD4ejxHGygK9hxsQQ3avWDESqk1OY4Wu3EYoycstzmxudN7zYj3jfj2s84eh8rGjUzKlmzzLl3aGn7nMIc/dF9bb5Exp8pRVDTUlXPVMsV9aDSH9tNF3mxVBQedA1A2HSe0oTFWiMALIIwu05hTtRVM/ST4FvBhRmnWWIdTYitE1WIeFUBO9JocQTLQGdZYQSrGEtTRp65ez9cP2kK7JKG5tDxtnPb4CpcRqdTzNWWEpYvukeaO30OjLzRb8plrLHya/VGPaSKvB7y7885/TTl9NBtfTxVFy9MS1JT0lRmZeORjQ2LWFUvGXsGnNyUzlz0cwAsLtHLHn1NOo5ff0lKG00Kw3/AEkP8ZP0yPJ9E3b9ErGngnLNPOkYPjSLhsxMsurmVMU15iIWq7kdGPUd4HneQBmcx1Y3yDDpqw/bT4FDe96LfuJa+/mYd+lzp+ZuruuBxprThrDbeLbfMoTBBqb0NmW5Lav2RmwLxwTMo0utYJukonNDpU0yiUyWR5GoBDtwpiIPdy7zjhWYIT0hDtGR7rTdsRatIJNrI55s2ENpQ/vTKMgxEuMFSzLWksuRJ306SJguyGp8qUBxgy16SP6mP6ubL2IseUZwydxWkqCRUchugs4iYpPE12LoSmhhiGY6ErIMrHaQY3vzKtdjBcYzqI6iE8oetAsQtTIdmEXKIBPl6PM+nUmcukYCGvAKcuAQm9hhlLMAawprL0ipU0aCXZE9F6Y/gO9DFpRqE8ooGEHMFvnjmLlFEqRKtJliABs8CTHE5E1GKeE8OH+aCLfsy7Eu2Zh8aBx0zFATXmsIMzshv5mZV1UEeYKDLMQnx6xG7tjxUuIquxL56wDMv098v5nX8fOfM/2UT5t+0b+V0SvJ4GjGS3BG/gslAzIph1hrQtZuh5lRFWUocgwqNn2kOT6Icv0w5/phXn24BSlFdQkCgNIttZGOVg44iYoxaMFzCTewhDobktN3FQuPY7pM7KMq5hwI6H1Tp/VNyfXED3ma1UCht8+sIhXbw4lOjdrEDwJDDAG5E4t4dZ52YAwXO5YXMHy+Tu/Cbv6p8YzVD6MK1nVT8pZZ7TH+OWDQ+RtAYCQmG3IKrwYMseJUmCDuAVNDLF7kuAsIKCylg2HOIvn0s5vBbXLYPpRiForDYOJhgaYEGsHkzYexGdE6vHWBgxqVfAIh9LMBKrNB/wAYAsPnBrl2KNqK6iiC1KwKZnaOhHSo1REWAEbxzWRfDynW+k3L6R50sI2Loyx2NiMhdC7QyHqJQFjBpecdZ60o2Srd6ppiNLsLGD06cQw0uYfhqfomK/jY/wCSxLKHlDap2TOdGCtlO30gg3KYo7kDZM/ZR1Z+cYWTRvSM0L2m3lzCH1ec9koKmEZ4/ZjtezK9PamVZeQlROjY2mFBS0wHQqGG4q0SV3ReExvWuXbJV6eCCZzL2oyn0R1opskwBKiTdWayoLRWBeYt0txPgOfFvdT3fh0TWjvPoJr8T3yMnh7WEHje1Zoe3gCO83/gT276eD6HwbJojpNWe9T3T6eGrxI6wnyeU9rmt2fSbx08f1U0p9t8P8vp4mcR1mjwm8+O4miOng+/8K92+s95NRPf/B+JxNTvNLu/WaI6zVGfM6eD7lPqfGOrwvZJ7P6Ju8B9VmnxaJpJ7zwF7bNfwNaavKbZvnvSfKcT6H6R08DSbJrk+D9kn0EY0w8O81p7lPYT3HwG0J9TxvX4ftGak0TVNLt4T2kdJomlnvv4w/bnh//aAAwDAQACAAMAAAAQfTefaSawxCUMmhkCFZlottdENJ+T+y3/AHpplN8tskgNZ4lEMkkkjsllKszwKSIb7bQZTaZyCJihUEr9Xqy8CTK3trRssuCaCSIW+T+/ll/tkTa//aCTSLVi7llti9llkMm20P8A8i097JLrKJJ9J9/vqkGnKJc3UDNVUIGko/vuZqJLPCuk2gdV0tt9ICL9v/8AtBtpppUsYSaSyjWb+62jIMgN+6ySySQ+feVdrqpptqyyWboAuCa08puhJx8bwUSyUdIJJpMbdq3727+TbZStpNJBEPwswaOZf1l5MpttJWyaSXITeSrdRLBpNMi2X3/AB2fiwpJpp7kb6WwuWWjqoN4tokPfq1wxezbZSNtJNNgNgIq2c2ZNNt5NZXTz0UkW7UooAbtNt2mTyPXIM2j6SmApp1oaB/f6a7S2U2/6fNtFNcWWSyX7/MwtpJNtoxoNIJNppJPg/wBkooYp323TqSzLbTYzIt+WrzYNE58jYDbRggWF252uV2lltnyza7Sa8tskl+3fXbCSSSQTbQQCbIXyS7trW3+ls+//AH0gEmmnCLJNh510Cdb8vLCC1RWm3lvlJt87/rJJNe10gcrpLLt9tNW2yw0wGUminRwc+9tPKNbv/wDf/blNJtppOLW2S5bT9pAmfd6+wAXQkNMJJ7Zvbe+SEWz5d5se7S6iW/f2R9pJNIsgJBuiDLf+/SQ+bb/b7i7JppJMvmWWavb6rYEBF/7iWS23+IwtkhpvDfbbu4SzzNpqB7zxWX/7WU90FbokAvu997X3aeS7/wD++XGzTZbaLMJEs0+e+n7aBIH31k9l1klkhACYJT+rX+28MsucaaQpexkltlkknthOTab4In1930pk3/z2+KwbYZAbDxJkls3H+2CQBBM8+wIsvuMThMoiTAbS5O380cmkeKTElm8sckRnttttLatmhgSYtlpIk/3XfY3zbJXNwJtl/wA8ff8A6XMskI//AOyz+7bkXsgBpMQCTab/AP8A96SWYN/95fa2Ryb1G6SxsgAiyyWWzSz77Nt7R5IJMKiGWe3ewmb77/5lEgvS/f8A6+3RsWm0JvgDKabx++/1vlsOKaWK/wD99v8A2QS2GqS2SX2WWNfTb9JRlJtlMwX67e3Vd7b77ffPBEFfff8A03sX3mf/ANvpKdkE0lnpvk5JpIGA36n7v9t/9adTbrbZ5Zqkk/f/APpNNpttiWT+3W+/P727/wC3qaCJGzVu3285A5jaW+31lhSJJPT4u9yvsoPTXSym3+/+2/cltskxq2/+30tliJSaTwEl9vnu3/z++/8Avp8wwCNk202n/nV9d/sE9dJQWwiWm13vv9f5RkkxQ7Fup99vJWlNFf8A/bab/wC+SSaacsl9v+2+2e+9vp+2tqTLBJ5SCS7S2v43+/8A9vb4aACUWGk+1d9LdbaG32kk82tbL7ttv9P/AOu6awp9ptjkyT7ffb763bbaf+eLNrIEnwppAIIzr1//AN93331g1kBAJAaX23XlskTSSbZTT7y/v328r+kzDlqeaaZCWFt3sy2bd5n/APt9Pbkv/iSeeSQUAi2ZnrU89vcv9tezQAUmnk9et/IKESESWQc/1ps8Et8k3uE332wUizLLJPP9v/bd/wD77fadPZNkDQcAgAgEFAYVpPv7ao3feQkikFF/oTPe2mEElkotvtp3pdvttbLNIJIBssGPzaey7b/R77JJf/8ArzTyoZFn9NIJJJILyXCH9V+2f3+38hgIBHz0f8ugMtLEUrIaeSTJTCTbSDYZKSQIlt+sh+umu1ydtrTX2aybbYj+ipsHLfgIWQLaFN5X1ib33v8AbAQhV/O+rZSSyJSTASz+CUwEgkQSGWgLCAVBbJl+0kumgmQAf0bhQmUAbfBvtsGPYAKPwSSeF8/t599r7DaSRU/5/wD2b+3+2UtoBK0qWlsgkkgAOQAzTTbbf5Z5IAgiPRWpABAkEGbeD7b7/wCvMPPQJIBID5f38+3/ANcRAEU/5ut5di+5vbRKTBSoZADTaAyQSBfZ99/9c3mGSW21XGgAADAYZdtRv/tv9vpNPt0ACACBPt9sut/9cCGknpZtv9+tfrffDNb75OKCIBZGTP5fknrvi0AAkwAQaWSSTJATZttmf/P+/vv9saHhrwSAB5t9t9+99cQGE3/sdNv/AL/P/wAuvf8A5NtZFgBpLb/1tt/3PBmAAiSCCWQflbtdZfvo+prp/wDPb/w7Y+2XokAA/b/77Vf+GBJB7pNJpr7V/PK/r/8A/wDbb7dJ/wDZbTbb4pZkgAAMEEkGyX7/AG2320mQ3e3v13+32s2G285JADv3r+38W9uAABIDSLTAO/8A94/lk/8Afb/b5bZqe/7feBskkEgEGm2UaT/b7f8Arad8H++//wDF/wD4nsp77E3EAkEheb/7r74w4AgAkEEf377X/W3y6fZv7Ta/bbbpNIAMkABcmEyG777b78rpe/8AgP2222+GB+C0b/325YBJAKTu/n/29sBJAJAIA386cYKvim1/++f+3yy+/M4AJJJWWMtt833yfjxie/8A98Gv4t/t9v8A7hY0ozb7rMkkgAbx763d7ckyhmFf1nfzDe03pNXb/wC3yZvH9aIAIIIE99D32X3/AHn/ALCb/bbVkEFTD27ff/EzutHT7fIUkkkAeff8y/sNoTzRl3gF/HhWyPggDX+drZD6kEgADLVLLbSbfNJSvfbf60LCpgEFVbpjbff9qIb5XT/bd/oEATq39fdFopNvygIkG06VoEKlRb/yAwklAD7bGz//AG3/ANv/AH2ffb/ySpUElIAEk0w0SBT2Fzv/AGSv+29cFwJ7CZVelLVhD4VfFo3Sq1zi3n2Pp0jYLgRx3/t+/wDtr1s5v9/t/r2FiACTsAASASAJQbt895v/ALZX7/7leRVXx2HknULxK8XYAupogG5GBqjcT6V7ONCeIeZYBve1e7f/AH/+6kIJpIK6OBBIAAAJJp/NtNm/3hYZQ959BJHFgQE+O1tHdmnsy01GDbl02sORYRJb47OEmd/++++v7f3285JJJBLa/wA5yQCSSAQCToEQP1Hngx7UDk2huqMQAm+aOCWUjp0b3AyB29vUiKdoRxExVvjvq+fYGGCKBEgAC2zXK9v9mDY2CQSCQZO4tkg7XVaRlYXV6dulzbOuTRgn18WRli99B22YeMMaFne3EekaohoPMaESn2CQTo++0vvt9/8A5uoAJR7vHQrjyNzoOwLaEwzKpl6uPdD/AJlwn25tTPALA8DkcOpOoRVN1NgcB9m6hhfe64JWW2X2/wD/AP8A323yBJeCxxPlmfCRCEdwPI4qNN/LonLpNsE7+9Q6CnWraa7t99szMdrrRmN02Nm2cLiJCkIXHW+196//AN9wjeat58mzXkaOdDUfmjHFiZaAd5jkyxAs5suy0CHnluNA5XjCm8pS8UeYIIzV9cy9RGilw3rycGNf9P1qaJ86R25gQRq/NBOPNa2PWIzirLOuWBfKtKECXQPsG8Q9kC7cUVTprQzkxIa94axATjhZdzYNodRamFLi8mq3axpF7Sl8EQPz/B7n+ZjLVfizfPBDvKyXDBFMRQljNwp5EwqIOEB3wvkb1LZceK+K5nz1cCVXq/Rv3mNg0z/dzppDAWwHzQl+JltXb8rDmEg24jWQXmc6oHTSeFb182KRLC7g5ABSjzAebAferO1p9e4BLtvyUPneKDlNiErrWU/MvpkVaRhB23qKGpfeXjYIC7gZ/eAc3QHhlBqjxLuD5n0OG94eD7iFFPRF7fiVyhulociq4Benld6q0RG06HdK9IokCk2r6bUl20Js2Tjy6QDEcdxkJqw06mH2NeUSdvfHBxr9h/bbSQEn2GSA/YYIpMZDjnlsQv8ASwadmjSKT1gsYY2ozEib31NGVUZEheWsnShwozhlq/8AAXNLDTJVnSEYUG9HT6q1FF5r6XXLoZIbd4cyvQc30D/6LNBmn5inysYPbADXCQnsrtN7hgtdPiH7NYLqyXyS9eFVnFrvjSwHO/CYLU//AKTVsF2n/hPuiUAFYS/+naLjRvCuPAM7pN3LEjt2+8z+pQiCu+lmVP8Auo4TGCx3t6qJNiv6iYak++ctHtO1TPMDX6sTyem8hotuh8s3ELzeiJ0a1m3SbzM/lBELMGb0YsJmXpRd+2tYkzfgF4UyfqeA8JRJcU5Qz1MjliqqSQfa8Yl1qr7Pq4chZPhmg/zSwPj5aatlBGYkLbugl5TJjVS+Pji3P+x3QPpsYdsX0dMD78es8NSMq+q4wmMs1fr9s7wRWQbIYNOVxDE4Dz1xwIokJfRpWVWnbkDS2KJMNHTrClJ4ZenspdjKE1gmSUyVpIsz2ilkgvdXpUqYRYnRkzYRNZcKMsQnl2sQKXPiZdUec53G2cT8jzB6ZqdbbHgjU0z1+xOUpc454D2pGMGm3QltqLpdJkIJLSAS8sGxLNcIjRLF8QEXaFdup1+2lPa05tOPZ90fL9B+V6M/FQ5HtEAfohS0dyb8iXcC5KDxa9z2GWtoU663SpY9BE6a+biYlTboz9UL1zXkvrOQx2HsGEBubrtiKcLxr5erkqndlSafPzf0lHsKJt1DNk2N7qtcewXyT2lQi0eAlM1yNQy9cplhGDZeuQusd88DYqdFwFYOoAfN7Xr3Y7nLEC9Ia1nccUTneXwaa+LUmPIE/wDwXNI9JHhFSqpJp2kgxSZT7PCXxyTIM8b2JzM6sr3pDjRbk7ZbZo2PLOqqBkGk9NsS6/RRI5v19UWWIuV7qlzY3Q6eZI+ofDjPO2lh2QmfKDNZ7gaszA2xJreKq9EguzT5qYowvnXU2phEccvEbEvdTB9+WK042zlneejH49LHh8XKTAOQFeJA2wxlx64HkOXhtnhPFMvUTmO1x+3CVzRsLF9gZPtdgSrZYXQS/wC29iPkoJab9tmJXpASUqn8LQVZxln8KL3xGdhsNB/sc6gcwzEMGS6zezCeQEPEVaA11Tn2Iu+uTHH86jrdTvDf8nh2hzKkU57xoLv49aFPCUCpGdDxwc0PGoVSPRiUDesLA/T9x7tFULok62LbtY8X9nFJou8tAgb1fKi8tTz2I9pKdtNLrFzsmaZv0zgnY9Jj9FApMmiH28vtrGfCmw1LsZP8bS09+6TOnFYJP/yZxD9DjmK7UiebaFWnDyL7gi3HXOV/lwaKAsnN6eCaJWSAe2oiI3JPqCBkEVJqlj0e0QT9QsS33tUlOj+/LeBW+AojTfAjpxbifcSJqUh1heerO9QvFYcmNkVVL3wKSvmhL8tE2knm2OStjgsnZ/oLgenzWSeoRF8mG/OPVC9JwnXa4HTADqeKB+oMYMxswqDrlkF+HiaRCt6GBbPwbyIoC/JbL9zAuPFPssh3RDjZvQ/WDZaLVN8LVL1tDcnkNy9OHruybyE2t8P7pmzH3F+arw/WsRY6UAzbnOxzC7cGcuNpOPLXPeD7ajAJna1ZuR1kI+pwWv59LCUOaE1N8/B3HuL8R45Tr72u63suqk0BjuLtjlUoIPCZrOU6lN5+IhHBuBXPSl+M4I9EUIoBwFz4zpxdsTzJzL41Hy4fiPT09xBqfqdEpD2gGlgRAf2Qu17TV0xCGkWU+aKm4p7ka4p/wgM6wY4bJJIbomx+Kqsw/RJxOdzXXEKHasu5cGQTU85ROHtmI6HEdFbrxyHKbKtL1ZZBzbLNAAaaD5eC76QQ+vPygOOB5GqC0djq0esNJffzLmUPpa3Qf7KrfNqQ8vEXdRpU+Dep8K9hgRBM+H/LNP8A6jJagb7z5VcSTBR8NtT2ApXdvuTJ638ZynH7T9HAb3+cKP13lEHJvNdvdGnZ9AjTwI0ak0ju99xCVpr1Tn8CqENHmnpqBTP+BnqSUvF8D2DUU/5YRDiaTDCoEvYE+enlbcBofEiilHQuNA495aw3PI8II8aHnjjt8uBR/EiWy1ZnZHHQV9Zyy03nhNDS+HUj5QVmiANMKX6w05llj6sh3O9IjQysv/iqzS1rAZ3FYrdXjZ2c04wJN4Vd+C9xpddCUQxhaVr8B5Qg/Wsw/PrsRA0IOKlCpl0LBqA18a9nv9EjgFTN0nQ4KRTxwIPblmvi1h2SfNvDjT3eLZcZlWBuzES8+LlcDQZEOATZeUtxlnX1sdvNYzlKroYbHCcB7mnDdV5CLpftxgeYo9CgDOG21mOH/wCndwuGcY7YaQhZwQOfVErR3UBnmMkKCci6tThYCy2eKceJQWUEKn+EDbJZjsSQn5B5YifLnvLnt+94+vHv/K6K97UNFqkv2levz3l3sGi/mAFle/RHYbINGNTTYpkjQv15WauN8qpmpZTZT3A2MSxMRQ9UBeHwkebxi9spd1F3JEINFY39vqgIoId6Dx2+tkl2SNBYXqxOmxAajYXa7wAcrpekvTqAG6rHbWw+thAUuBDoaPAwozwjMe0v8q+YFGBo2++HAzyQ/mbDBbFLU+LnbAFXkiC38jF7aAdhf/WcK/jinGBkub6g778/MJo5RKceodQKCbwTT8Vl0zI2r5yyAk5IiS21hX5QeweR/oJJHufg21A1lXm7qDTL2gLtIH454B+epATRAjvdNxXwacLIglHeAzfSVWyoZ61sdy6lGIMP8dawpYk7qHYGi4nYP6EyXNhrTgUjSQOfiuq93/rL9+dsfwcWFPTUU+LEmsL12CjX2plEJSmi7WEVq8AVpGIeacTrbvfyQTmluIJPZ/i1bxHxFcUlyy9zrFW72JEPgd+Idx1Qw6c7J9eiwvPxIM6i8jOoOKNQ8PpfYAR7LfhYK3ySWH+XD1VzTJVl1kkvFqz8nwjaPo2TKiATfic7xZlSo8RtAB9Tuf1HbT9Z0s4BSW6A4r7eYxPU2Icb6V6a/DgJB2j9ZGU/Dv8A0DrAlznFoOwwxj+Kg/VCswRtl1t761YrZ/gTc5J8fDRjc3KgDAobeRs48RJ2NvXSQlOumTwEJX4J5NZtREHW02Ldy9HWnPsdYvFx4OKL1iNnRykeVGLhEBrjMNLSqk3nI9KFtVcvmaNb8T13n6E+Pk8QIoVwLoyIzdqplKfR8Eii6CedY5sxjDGr3Sm3jPAd9C6Xw2P31rq31EQ8rMKn+XFMkjXJn4bZzA79iO+jgs5Zq7VMx/cs5XpPisvkEFqc3mRUadoeH8IWEB9cjJYMIAyFz07CHw6AL02tJ4GJ8Ws7JmwlJWyjpKVG7F5NMPA1kk8WJhsyMfMkhndvb6TH1tNFdp+APsXPttVHPnUT/wBNdn4YeI2Ke8Ex/wDl0NUB2fli/wAx7uCaBp6IgEOhn/UEMN0OByf9u+EwEw3hrp3MuqqVZst2gBFWYxbSORND2oGTftkUo7QUKFHYIOUWsPNoBwFKAkNFsgHzATI8u/t4XUQ1z0UAry5OoBitasvpwcF+m0KLZSLD96aaQm/n8jU4UM5o/wD/xAAqEQADAAIBAwMEAgMBAQAAAAAAAREhMUEQUWEgcZEwgaGxQNHh8PHBUP/aAAgBAwEBPxBF8nnHmHmHmHmHmHmD7g8g8g8g8g8g8gXcHkD7g8g8g8g8gfdHnHnfJ5x5w+++Tzvk875POPOPO+Tzvk875PO+Tyvk8o875H33yecececed8nnfJ53yed8nnfJ53yeZ8nnfJ53yed8nn/J5vyeb8nm/Iu6+R9x8nn/ACef8nm/J5nyeZ8nkfJ5PyeT8nk/J5Pyeb8nk/J5vyeT8j7n5PJ+Tyfk8n5PJ+Tyfk8n5PJ+Tyfk8n5PJ+Tyfkfc/J5PyLufk8n5PJ+Tyfk8n5PJ+Tyfk8n5PJ+Tyfk8n5PJ+Tyfk8n5PJ+Rdz8nk/J5PyeT8nm/J5vyeT8nk/J5Hyef8nn/ACeT8nlfJ53yLvvk8z5PO+Tzvk8z5F33yLvvk875PO+Tzvk875PO+Tzvk875PO+Tzvk875PK+Tzvk8r5PO+Tzvk875PK+Tzvk875PO+Tzvk848o8r5PI+TyBdweUeQeQYNjzDzBd4eYececec2+/0H6Z6H656J6ITpPoT1TrCfTfqfpg/osX0kNdH65eiJ6F6YT1oZPpLo/qr08CKbffo+r9E+gx+uEIQfqZB+hL1P1z6T+mhk6P6WusIQX0YQhP4M6Lov53Aum339L9MJ6F0g0Qn8OeiE9LIQnohOiJ6YT6MJ6GLo/VfRRfQn0F9KD6rovXB/w16V12+p/RnR+qE+jCE+lCEJ62vVCfwn1fWeidZ9CfQnohB9H0gukILojjrCEL6J9JDF149C6rpt9b9U6oapPpPpPoz6UJ9TPrhCE+qn/OhOjET6D9S+tTPrXVdNvv1nonR+prpwPpOsIT1whPoQf0X6H/AA2In0F9N/wOfrL0snXn+AvoUpt9/pPrOqDRfThPU+j/AIcJ9ZemdITpBdV9BIfTYvqrpPqr60F9NelenaP6TROkMdInRk+k/rv6F6Ifonofphs19R9cl6wnXZOi9bF/BRBfVnrXSelehehdNnpn1D9D9CJ6Z62Qhr0z1snR/ShCdJ6162idIT60J0X116F9CfUvqXpXq2+ldH6J6KIb0z0z1T68J630nof1p6p9KEIY6QgietfSXVfTn8O/SptL6J0hCdYQSr6F9EzPSeuE9M6z1z0sQxD6wnogxfVfonSeqCX8VfSz1n0IQ0bF9BL0IfoRg2/VSonRCDJ/KhCemE+g/pZJ0g+kJ6X/AAl6J9NeqdIQS+g+s9MJ616b6tvSfTWBGxL0kh+meiE9fBPov1T15/gIhPTP4Guk+jCdN/QnpvWdEP8AjL07er+hOuvQNT1NdX6p0n8F+mep/wACdJ9VfxdeqeqE9M/jr07euxE9WxC6pjyP6T9UL1hPXPW/pv0T0If0Z9GD6L6UL1hCfwJ9WfTf09v10r0IhJ9KDXrXXP0YT1P0wnoZCdJ6mus9c6Qnon/zl0ZOkH6UMnpvp2l+sl0TZt9SE+pPoP1Qn8Z9V9KeldH0XSi+nCeqmyfw30hCfVTL0IvonSdUI8i0Lz6J9J9Z9GEJ/Bf8mdJ6dk60hOi+okX0wwT6i+gydF9fZ6oQnSCITpeiwNj39B/QfSfRvrfpfqf0NEIT1vous+gvrTrCfQX0J0hCfVX1ETpu/gLomB/SnSE9N+lCel+p+t+iCN9L9Bi/hT1rpCdYT0rrPUv5+Td9dGxENVDUGv4kNfQa9b9M+s/oLrCCIP6MJ6oMvroxD9U6TpPXP4fHWE67ukJ0hOkIT0oTyUeUbDIb6Y6wfpa/g8E9MH6H659Fk6z1ci+hCehdX/DX1KP60J0npz13fTnpQhCet+iemE9TM/XfonSdJ6IT1P0wn0IT6jF650gv4PHonRdZ0hr+Du+pPSmJjyNfwp9Gep+qfXhPqz/5E9C6r0T+Nu+uzPWDX1Z65/EhCE9c6z0zo/QvoT+BCE+hPTPROkF/Chj0r17us+uujGhohCE+hPoz6E9E+jCE/gQn0n6J6YQn1IT1z+HCEIT0P6C6b+i6TpCE+midNvTOk/mQn8CdZ/Ag+i9EJ9GE6zovTg4+jfqL6667ui/gp0mBjX1n0RCet+mE9cIQhCE6QnqnRdIPpPTP4c9M9SGhfxIT+Cuu76b9aFjrOhr1z6b9b9U9E+tPoroujF0n1J0hOi+mvQvoL6K+pCemelcvqwhBekhHH0ifTfpf8ioe0x8DGtiRTCGmlR8KzJJjQtooWDWYJj2J2mYF6IT1wn1p0n0WLq/oL1onVj+nDcTpP4NExPpDtEJ9Br6UIT07J9GEMGB9HtMaeSmhopDlW4V1vA3XENzEKIZ1i0vhGShZZGkPQ8qhpZLYncaYn3Y9Z9ElTwEwTORI9eqfSnohPqIvohCC6T6e+rF9Pd9KfSpSibF6DIT1b6NfShPTCEINejaBHmjXhDboNbY+eVLCyTkJnjQqUSbdDZoMKZuh7hyLCMm2Nt02ISr2ENFvwNXIqw9mdDDyjAZWhtt7Kwl5QW4LkQuZQXKE7T9fHon1Ia6T+DCC+pCEJ13fSRCfSQhDyNR+l9J68DQifSfSpGwYlyIaRpA2sh7jbIlsvYYWxW8FRzsNMEU8h8EKN7G2BKIh5zgfcyBuI0o2Qsoxgo9nceUJvBjpCjDHyRkFZCp7RhrJUKhvRWtmGZ5QkbHKHLSEvIXchoAmnp+lemEITqv4CIQn0p0hBevd9Hn0wnSE9CNBMafQwf0J0ZPQ2l0Q5ajQGOEjRBsiprI234Kl5MvA49zLRdhdGDkZWmEJJpWgiQoEQbMEJEcTbEiEVFyJJKIZIYIXIeoxKoZghqM5nA41CLocajFoDj2VvocFfsE0tMOgytEN5MrTIezK0xppoV4Y2+UJJ6E9BgEEnyMDbGmC1H0Rj0z6S9U+rCEZCfRTL+IuiF0aF9T6MS+g2l0Q5aieZmkQ20D222TtngqRhwZaUGi2F2QvkQwhTbMZjejAkyM8BJt5YlYQmyDaRn2CiUQxsEiCkojWWyjew6NWl0emaRjU+4pWAt6C+HsaSRnC9FRHkEug+SwKcBpMr8ipImhJpnciltGWjApvBGtDfYKPYrW0X2Eb1ks2oJgjt0RwDOjOUNML6kQnSdIcEIT6qH9XYQn8VCUSE6a9bINpGnDlqPkDgA2UD2xnmYsppHGRDSmWzDZT0JdsTTCQk28GwzPQp9BvgQkyEpxKvoKkivEaAQE2XRV8wpMDc2bDXAjWbJCKW+zox8OmIExx4Nr0dY2QUceBvllCaYhurYpc2GqoyPIKxpPIm9hUmjAY6EQwK2x80ytbKxHwdjQknpkQt2oR8MqbVMIj4J3QtSDRBK2qIeA2jhpAlMPrP4cJ9OCXTZ1hCfwksiKLRqdJ0vQTnqcqZpER/SDkmNdsXAVtIa7ipoZeBpLYqWplvBNgr0I230KehmNAbNIdzyNNi+BCRCcOSeAJJaQlYKeejhTJDOxRrZSwozl1yLBRP2F0wSwVDeBnsUSiJHSSraFCjZTQKsorZnJaE7oaiMuzQndCIXZlCzyOtdATTPIWhUHAbNldCNaY2W0QI1plrQw9GGmVyiaGYaG3yjD0zBYL3RG0xYCq8DDKclejOEa6EW4Knz0hCCH0npn0Z1gkTpDZ64TpCfUSgskI0gY60T5BrgHzoPvf3GkE1wI3Jjt0XBB08sw2zwDTcwiZbPAOtsiZZhrJltkTY11kRt4Egao7mBZCEovgEi0NEyXThCSWhtLLKxwQjFDY2cELEUe3yC1i6RxsKSFRClsSCjhUwUvREfTgxbCYyYuGXo03vHSsaeQSJjo2y6k22GLGDMj5opBZyO8oveCTQh5RU8iVuDR5ImnSORo8kTTFO10KWmQ2hNiuGVNlNonZmBVyhJcEF7omwx0xaLfz0YntJiUG9uGhC1GMXonrX09n1Ic+qpbNoh3Id2DXAMdplnsy0i+5NjO1CtyNGxIJvgh7ZpIthDTe30KYXIzYGmkXmhG2xouS6BJyphDR4yJsCSWhHIviQshDjLKNKdeWVmotibJyiEq2J+BfsSSURBjfIQFZBRHtsvR4/HV2vcJEOiEjfv0jEivrJCAg84No+rFlCpUyVE2AQ1cQmjKEM+w4dFpxC0avAvcEjGj4MEMdoqaHReCiUNXwRHgcbQozwKgkeyNka5KW0Y0I1plIh7InpmVplcroJeTI1yQlGGkK3M9CM7TRoAtZlT16J9XZ9VtD2kOWpyZj1hDu4NgZbZhhFfCI22RNsngr+DLY7op6MhDbGi0yvgiexeQt4GW3BIY/Itoh7FWg7CdtBIRsxsxnlqKLTEMNifJELQKu4+GbOR6Y4YhK2PtK7mlPuI2Ez34GCoq+UVp0wJXeBTohKixZMGCG0jEKVDqBTAtQhqmBmTowNUaYfVrlCHgo0nwRhNM+wh5EwJplXYbIKcIVCJ8GGsiTTQ49oaPQ3wUSyJ7RS0VsiHhEPgw0Y7Qk6CaGO1DApaKnBnsdETTKm0Q9ngKCltHIPBlQtbXQiY2WharEAhtXojaOGiCaen6UTpB9NnraLbNv0I5ExjgO1DbDE3Ya+CVsTIkMaFNiGyeBX0oU9sc4FPSM+IZjHaZ6RH8CkY09B7TF2COzjIs62JcOiXCoJ/ISa0coujAoecsyI22TbhCdTIjDk5SLsKMIyiiLLE7V/t0zuj04tjE+Qz3M9zQHAM9GbwmJFKZ7me5gIXuXyXybzPuZ7n3MHPufceeRo2L5PuNJ4onMMvk+4y+SruY7jS2mJrlmO5juNLaYu4x3MDAk5MDSeBxsJBgbNiTWmTzgqZsCPRkhM0RtojWiVoJHoYRrTEiWAmaKZMi70JhQSaE+6E2wNcCNaE3KK2xpcEa0Vyim0UyiPgrXB3kRtIoj7GhI0zShLeRnAZ3joBazL26QjNw0W2bcc1RaLQEjZhgNO2LtEm1gXeGjbJimhJvYi7YkaGNGW2Q2NPJTeEZbYhaOS3pEuxHJ3A7whLtiSNpyO9Ije2JJob2Y6wEyZiekQJ4WTkY6JEPdDuYX5NB0J6y6VEaNFQ8hleDuaRGOxhwPR0hV2Kuw+OxCKuxUNoSSMdujaEmzHYjsSG7Z9uk8Cw3T7H2Hh0+x9j7CVmydUZ7F8D9i9NDVFUJsd7DVWhXQVaMjV2iNaNo+jV2Yui1sTuiUwzgVNop0d6FPkS8memLp0c7QndMaMiaZHgyHyFrTKpfPRfDJ3DRtFWFHHIkaZV2eRDEyWH01yRhdrInJlbMCVFVyacbBiXtHsHkNGx7RmZIqmWhlxCeaN8RD0hv0iPkEuIk8ItoJNs8FFxBs9MNnyKuBHCGzShT2KLSGi2U9IjbElwHG0S9KjfiEkuCuwlbQnpUFlhRNrCQ3W0VppsFdiPAIw5PtL8idUV9h8xoL9x6dyZ7CtcEMLZbfgZHRslSDGhIwj2GRmkMDF5DbWRm8mTJWVgKrBkrG3C0isyVjqFFZkqCbIyZHWWFFZX3EZRkz3MjbgyzJkyjJnuR9Cq2Tsz3jvY32F4IQxymVgTT56NXsiadPLBvkdbMNjAU5E8kkTT6Sj0xozHTIj7nEzD5JFLTMNiYUI4ZhojkTYgk5K1voRjsMjXJfB3ShHDIVLaE2IEqK5f7KLCIxtnoPEU0iu2LZBxg4yIyPNUsaPFFtIrs4CJMjZ6RW8HnkrWkQOMh7TFwIbDfSL4DzyZ0htrYsBDnDiLo5bOKLbrUysHcaHI1vwhOpkyhu3My8noqjIzJmnocMyZZ35WQyR9zPcbaEw0+5H3MmWJObI+5GOiTIzPcjEmxGlgjJ5MmgjKIQ2hCeSu4+4kEiEMPBlYZBonY36NExRK6J0nZiZfPRq7I0JpkRgaGVvImmYMDXacE2w2QwNha0zDQVEQzcB0S6QVjTD4iNayLiCbZQ05LTMo4mKhhHDK1tC5Cg0Ilpla2d4rFDWmYCXkTYx2J+6/2U0h0U2LZBwU0hn8HcyZQ3QtJD0UXeVrQ5E/SE35I7DaDctpDZtiU0UQ5OBgp5akeiscaEvARdeTKwVOSiJ0vPEcBnuH5GlaybHDhGe57jWTrJshPgmTuGmuRqwss2HE3cz3M9xiwmJ7WZ7me5nuNsnJGR9yPuZ2S8ldyPuRiWaJeSeSeSeRq7EsdEPcNYCRPJCDxgSIQaGqousEj8+kITlGPcSEImLDx0SbIRCi0SkREQiJBURCSGjI1rIoyIwNGJJ5FofTA2E0OiXlQwY6BHo6KHgJmiCxGtMx2hNjHcbCNaZS2hM6KEmmVrjoYZQw0ytbQl5K3RneYRXL/ZiVwhtymxRpDg8VRttFtijSIDYrcQbNiCwijAXAht5CbRFDnZxkc4LgXQ2WzgDlCKJFFTY2biUeywQxCCiiLLOQhw3RgM3ZgzhHFJ0G2stiftnCEn3J3DvcbbQmXJH3I+5H3MlEZnuR9yPVH4I+5H3I+40+5HIRkZH3Gn3EqhLyV3I+5H3Hh5Yl5J5PcTyaEsE8nuGiR1DS2JQhCR1CbIhCE7Ha9kmGTqJ3DHBBmJNEWhMIIJEhsQQQxINllFXOBJMgaPg7ka0FRBA1eUTgomcEDThDBDQkWgkxA0fBS0VraEwwNDHREJW0VPQ0n0o1yUtoTiLpY6Z5hdvd/sXYJ6VNIuxiScGHA1WzLQp4JyVEi4GiGg9ZQjDLRC8RSdZb06RI0iu3Q6wieAQnWqz2FdhK3A4orLMTaRIrsV2IOJVjXhCJYkUuCuwzYm4G1KyHBXYvsPKIq0V2KKxsl0VUZGxRXyZMlFY2x1YWzJWVlYm26+ivoodHdIVMmTJXIqZ6KzI7T3FfcyZ7m8MVM9zJkTJ4FoZM9VDkGzRmTPRNojLoS6JCHVyZMlE2PJkjJ5Mtka5PcS8kEiSBUQyGrHOmN7EMEJ5GU9OmGkFwDEs8Rrgok5wSkvQvhmG0WhJcDZwRtEtF5I8BCK5f7M94IuXRJIcE8FPQrYJOYVFQhF1YIewkmiohZY1elFKtwSyoqNgzgvuJe9El4PIR3OeHrYGcbrPIR3PMKWMmTbnsRRdDyDVHCEzL1lRHQkbMTQnpWGuiqkkk9Lk6JJJGonFZBJJI1G4SZCJ6YIeDb0X2dBeB7D2D8OjLWOD2HsPYV9i+BcQUrL0Y2sG5oy9KWirsDGyUyUpZQk7THdhNlYmVijMorMsr7FYsmTJkyZKVlZWPOyO4KK4KZljd7RGtEtlvRXTLJthngx2J1YZkaux9mCL5E23gZPkjGhMnUxpNFIJt5TIyBf3X+yEsjRo7AXvCRwSNA3qhs4gk5IaRKGi2PyBcKCVbyJexHYQjJMmR5wZKERBEyJuZM5qI14gaMiRVMn0tBEiEIhqwsiY4lgg0OD7BLl9YjAyInoSo3RehLnobr9KVZa6/Stpi7+jXQselOMXoZHOhqqM9WLWNCjOilhekcZI2loU6waY0HKuheuy8GXoYKb0a6Jox0wa2VMwNoaRYLoZcmDHAm09iohCfQY5K1oSCe5BByoa0MUaEvpQJuJFkeRF/df7L20JJpE7RtNlcIb1YL5yYaR4DgHOC6lCmchaHTDsGhPWi6tRIRKD6bZbaE7jTZPsJCJIaMLXiIPYx5TfYTpETqGojzgWgQzvJ3DhbGexH3I+5O4j7ka5Es1sbPkruW+Rv3L7lvnA84Wiu5H3I+5H3EzcTNCruR9yu5H3GvJMPLITyJE8mHImwvI9whBKCSqpM9HvGiIfITZck6kGhscohOsENcA6RkIREQ7DglnUhCEGNgTNWGRqEERExKOoqBzngiIIiFqjIhJQgSD7XQ0Rgi6Y7dJNCa5QqI7ERA0eh8AqPt1SJI8ErCCbaEk+hBGjDYjsojXT7E/ff7GmTGj0pdjhkryRcERjk2BV4FcuaApRqssd4zEjnPYz0yYKio37HoYvItj1iUwNlG0tidLWbLiIiMFIGiOHR7oPpUNoyRCXLKulKU9yiffpSoST9h1haKVFLBoJOz2/wBCG4UbKJiQ6NlI6IGE9+4iopSluitsoo2MUtI6paE3yNlLeibapDzCwydh4BPwkR2jwDktZ4MkbHiPEJ2hDDRTYN3nlwNeWx4DwFdIoU8L9zPCpjswRiTZVVLAkmUONwYmqpDXloosaVSwdgbJWi1A2IIJN6MqkorSlrlFcopONoruhO3KhjG0LuIoauxPKK7optoansXaxNZRvLUKCVIbcK0Y1ErpjVLRIzkIapUh7i3vL/Y2bCo2LsNG2cCZbWEdgW5NIsHnOQzyDXmD4zvEJ2YGx4wNJtopzkjbsPOUVylnWhtujq5MnIaulBt3GuNEpD2X3GptkNUpKtQbSUw5PB9y1yNlyIsmWNJpTA62KhmUOinoTJWRuwwTml1bwOzGInkSeCHoNDZ+wxFeNFRFF0sgv+D+xsV9KWvC/ZR0eTXVhCzYH+nV4a26N56LmVISlFORMhsUGWXyZK0Z8Wow1SFFD1WVyJht3EL3o5S4KcjvcgJKMXuG3NnexZQyDn9ldxOJpje6WxOmRyJtoYuhqmCnl5QkLDqFpMNHlC9w7dGbVCmDMhGlHMgjK0NsGplkpgOBwJpiq0M2ov2CRMCumNPJCYNPgbWsTLyJMDYk1ZQtDwNHlDE6mIZCbNHGyJfAaPQ0LFaMAzjC1GYaQa+Bo2OYqYx9Fdj7swg2oWQBZCGukpyHDldPqiltXFpjThRrcgjk2A8dRM1c0ohrJNmEJqEoa0cjEgSPtoWQNoqxuDUhJDaRlhQXky0REtGypE7jfHTao2kxsbrrKhLFehs+jGhFEMyFPskaJYXSN4FNff8AoZZ0SqIQoukeyGmtoZEu/wCh9OOlSMGuzpkjTY2K1BkbLSKbwiOwTGDPKKdxTL0WhmyPcpbMrgaOiVBV6QlEwPTx+DOcNMokihIsMj7CTtEi53+xsjQsZ1Q6RO6I+xQtKDH+EYzA5EJmnJBxoo0GwNMBtVgSbFnDGjWTPInORaNANNOPA2I1k08jmTY2mdhr2hMm1hjT39Gm0o33jJt0an4GQEuEEoJatZHwCOqhMZDn4GFTAm3SOEHGxX0YTURw0I7J/YeUajFJW1Whtp4Bjz8sTNTEvGxEO4OQQ6MBNryVsxonUd4OZBtVsk4vgiMhjcMIaCjCZTGRxNuHsx41ml5O4PckpaZ3IrdRayFTI2Jy5PshE1glwI1yU2cldYENh6VheRxJWuSGRyUrXIsENOWYCo0+msPLrIZSMAM9mNI7ZSE20sou5WYge2DQkSbJvNZpYa0ZG02NkbeijcHD1oRXn9OlZbWlyZWuh0f4WR5bfSvuJroaGWUx4kUTY7ag2VyN9Pxcstc5KyC2M2lawNsYtU0yyBFaeCNt2I0EPYSv/Tu1uhOVMTbzyinsOajlAQgtPABbyc9OYAkrjsJ8MWNCHka6JmkZhXPcwB0RBaZGsb6YG1FVauw02KQ1ODnEjz0T2DFCoSz/AGGQ0UaNaG0QmmSmnZpEfgZxlHKWRDLUdaIVcGTEUeUbcgke8j7UV3IeuX+xZjk2BhkNN7ZgbLdDbOELNCFobsVyUURRJuBV1/sN4UMarwiNP3Y22rU2NmhY7jrOX0HuaeORoUxXVuGQxFKB0Gq5DZuqrRCcnsajXGF3FHLyx5db6M5wx4CHwowi1wbeekuBKZyeB1cHMNjm2ut/gspRJsSESwZ04L0WGffBoY9FQ22yNbXXYWFuh1OluoUtrotYTozY5uDqTaIZaKmOsvyNRxjEm9Gcb5MTWy08jNrlF6Kro7Rs7RMoZvUIT5UUZdUIaCYmaUqi4iYN9ZRejpYBxa9yJNLuR2QkvI226SsdXD3HGMP8CsiyLGCGqXlH0gtmnkamU4rZRFGry46sPorwLF08kJ01rmKTiwc7UvDKhHuROq9BJQyRyUI1p0nkgvIuZ3p96R/sqoRfcS6agm3iGa2JtiUTLWQpafcexvJ9wnk1MhUZE8UZy8GcDI2p5GrZ5CN5kIMLnL7iuwQgobKbrIE8oSwWoILJ5Yxid8kFbbG3gNkNHtFELdmnsgxgY0TpmasfitFZVyJdJjuMjBrRZfTL2i0cA2ntCkI9jXFvJGtj2RxkdgeClyQ9ofqoyCHnkiSyWLAtnMZq+RI5KuUJiJw2nRhFaUQkE1EfcTa0XuhJ3lwSKjMcFfAsuIawTaWxvuqR91Gynpwq7DZkljmcGI2NwJ9yOwyjJkJ4Q2e2JzJXIk2mJ2sjOrQyyGKdIewz2GYKyPud0aWDzr+w24wNvZk7D3Wo8rK5JCdlG5RnscSwNN5b6H+NFAtmBT7kUsppuUIuPA230fVE3Mc0oWdqmISjGysDz0ZtSMckKhZj9hppxSYiPuPYMdMp1GKeV5H8oyjVRC2Xcg8snSGyYE5q9h0oAnOR3HdN4EkunyL/AGN0qGV8DnasblFgauWWaKSiS5GPBEJcmIf5QGVYwi9ORoIWCd2PQtwNjoSIoxCHCeRrHkyOf7DsWInLKUZrolMfuOBkcAonkY3oYk2iQqTu7lgkJsXs8IIMvYUl7aG23WNwc/xlepyKqb7HIhjHIUhQe3dcLcZE1tz0bK9waAQxYaZQ31UqYyTCyQg8X3fQmT+0JSLyKDQ2PQ/2NNmnx1pHDY2cEVE9PZptPXVOOoUnMXcImNKFpx8rrBpsRyY7jkGaYZXX7DTadEGlBfPJ4iJnuRh8jM7XSEMesoS10HLGR5hDoa2TomytDCRUNe/YYrVwWYwx7xm+jGkYsBYzYTqJTwFF0lVoLEskJeBjU1oiPyX+ysuB9hztndIkWFvQIZ2Ja1B0hLAg63WG0tFPYTvZXWjKYEhSjsVhDTYbgxZ0TuJcKhLHghVwx+Snyp5DKLmHbUehQaRDzKvsO5sIjJqacZRrxCLH5jeBS2CBWxmI72o6hsWnwjN6xvtsZU3HY7wHgGN9rJRsBRzRFCSbSZbKDtGpvu/Rmxgaui+Q9hK9gi9xEcQhvuJbE9xp7IbhpRJ6ES2RXEFjLwd1Iy2GmtoUXuExO8j94Y0qmLJOjQl2itYZjL9xK6Eiy8LKgxUKThjarTky2pPwY1gMwRyl9hOTEQvMZ1ZZixqMY7EKR/dXS5XhHEyyDqcOSQ1S+Rui4NE2Lv2NxoWdDlXE3E+SKMZLViqP9mPKaF5Yv8CNozQIm58HYwf1MxrBBnSiEYgqsouYxMx62RuUWF4Hz2GcMo0cqjSeGbYtIllocCNsDEhxl5GtlDB8DTBOuDJMsa3En7M2tlYrlp/sY1hBB3BEiZLyjmwr+hL/AIiKEMm1JERlaJeGhzoJXCsziKSA36IMSNC4ijEvGMtFFjiCgGCGJ1h5KuA8O1icWx5oJSLY0og0S3kU/VIRnXewxH9hNHsaBDTqKXcIr8BogiD/AMIRZj6OmnUPQlGspkY4GxtOjmF6aEJmwMlbHYVH4h9mOln7CbODYIWgxNVVklI4VvfRMmdoRrpTIioGekoNvYZJCp/r9FCUQn0xjjD/AGMTenRodZHupN8gngXfkdE4D3CDGPAryD05BcA0uzGmeRttWyQgm2oVlRijJMB7UaiPD/JkhDKdRFyoqKZPgXEpPa+Akp0ZB/3FtGfPsN2IzZo8CSINDRtRMJOmC2W7jG7QkusGNMmCNQ7pfZDqLN34GuMrpCCk193+xx0WnkMlWlY1XQQjg60EqyNzoop4IWGlZl2wSSNKx5Fg22UclwRKx+434BxEh72QjhDYyLSibQhtEV35LijbrNDYzt4P4yHhC428eDCHnoIk6qfgDWi0tDUwjOaBkl4G+AXVD4KGLoJNSciRKGd3CV65naM0rbNdCW7yabqyxN4FiROmTG5K7GdF6a0ZIYxlEr2KYujqibMqXn99H08IHReGanTF56aELxPfoQg7+C+7I1D2QGhb8i9GtDnKiZQ5vA7FfrfYaaca6womIIIZtIJ9T7dx7NvRnJMU7TYI2Na4OVhmwXRoYw1ywJSGSFNiWMt5WvRBKMbtkSM3v4HiGab4Iz5F/sdPAipDVBRl9ApqJUNwdDYjaZCGm21/sJguSqMnkwhspoA1kojNCS5sZc0huyoSWxxobok2gXlk+xbEv/gpnOcJLSfopKx4Q30UlwjMNIuEi7s75Z5SNGrcY33QxjW8LZ4SjCrl9ihaeCFSYSKwyhZrjTTj6JnSDpFpWxK6EqmVsVW6xjQVkWCEr0nR4OTFhGecEIimiQzBJO4jBPuNSqyum40N4RE/8C07GhsBNJuS0XJgxmXAtUGqlGZcF7hinrkuEK+4TsmNNYaF9zldH2NhvsN9JETUYRcFmxhJF+Apmtj4cPo3APCWWJWcRZbE00ZGPMgzkI+UKEzQxqkQ1xSeSOO9LLjD7j+J5QpJtw+PuP6AldGx8BiRYQ/i0T2xXWomlq7ocuxMvRHoPQV9x1uvZj9obmWx77IwiffoumCuCNJfuZ2zEPRTF/YmvGOYgmn05Gl/4DGMELAmTrID50q/2PtVmEaFeRUOMnkjBWozbiEuhEMTyaUe1sRc5R2h91lE0Qp7RqXF+xrYyDMA22rIJvJHiGNQwiERuYx/qHKLCJA28mJC1RcGGNW0LAzmy78I2S9JbyyGLBeUd7nt0cmTCHKix0x0f6B/4LJwJpCojJr+xwZeBi8rK1rKsNl/rGLykosaIP2KEs0NmNaWBcOWMeWUcs2n9jlnb3EM80Xsn+CjfIpSeI6Uw6bsY2ml/vyI4T/fkQzQeDgyzlEt+X+Bj1jEJomHv7FlP/wQ1YeUKlmyhFSYYhKfMzz0lll/wUxv/BzmFqWiWHewluXsYnSIhobAJCP9CEMb0ITrw+4wvkrmT7jbeidGAJM4Y5sENbmmaFjmal2NYQj5IRDGsLwxYyR5Q9X4T8sUU6edH2a7E6NCqdRiQn2IS/hN7YxcRZ7jr8hCDRoaW0VLexqjnh7MSXJF0MRDeDyyN5YgkjCGzIjt2GIkkFFyiajZyIqBtLqtqgiFEK68vuMWrWNMsSpDQ2NUjrF26NVtZCCsMeAgkYQ3RMzYRsG4JgwL7KETkTliVdJB46EMlJ+UMatjuAQ0if2WX9jLMS6sTwls33C6Uy5hORfsZsOfcx60idVSv4RmMYXVocAZNmlBdVqryPfRmbY3J/SIlP0LHRjtVbWxY6MwdMJ/8Ftf8Pa2I3EMUk8l6ccYh4G8sjQ8pbEjQIQg0OlwJWr9iALloeo+TKPHoaUgngv9iiR6EPw9hDHAtLYu3og0YDJFswjAaTO5DJV6INDytBwos7HsRTUq8jQxrHTD0To0xDlV5P1APJog3onSIT99/skG4MNjfAnooWcDVIs/YeZEUiNDLoewJ+f8BBFCv/ww+CJckNDYxM0QiayFat4ErP8AwIXOykCQkNjIoUmxcMs7zkLb/IxGlciRobEm6SDQLLGZsPUuBoAtc/syIS6MfYaKbexaH57ROX50Ss/TMvsRM5EujPdGRMjwYSfIuCfgqsfgyyX/AILqn5D89NuIWx/4xJP6Qrsn4RE32FGMZrBYyJ0awWyNew7/ANhGTa9iTIuRqxhlp5XVrkdkcRZKv9CSf5I0mykqUcp8CU+N9YNZHqq3wJCp/koH7HUqsGPWo+ZCJ0RCk+4aibWJVqf5OAWNpWBFqfYdWH6Ghu8Eo+54Mks/JTbTxkeBo9wXSDQ0Jvt/BCSrl5GxTXajaL5RhvwWOsPrCHsOVb15GnERAxO0owVZ6R0vdf7HJlhEX4BPj2BJPEeMRaW1CrKdEJBqhuy14H3SeCIz7wSuf4GYEQmWMkRNiJDA2NiZkkrRAtCB2CLPHwY1aKraiCjKINwbGMCxnQ5vDFBFX/4PaLQlrg/I3z2ujdG1wIs2Gr2MWjc9hV6/cc7f5GPLgSJ+QZ7BjEVoWh7thHAMx6LSGTFPyUSPlmVcAkw27/2PYx5JAe7WjJxCStmckt9xk5r8kV/kbewaLw/2MedGl0ZqRhv3HNP/AMUXH+BI04G4MOE2Yf4YjadHOPuijk0IstCGw41oVzn4GPj8IZ66lwMBXWmJvuP067m/b+xjQ9ODGqr+B2yf9FFGNEyYPsZ2pjbvt0SbRMj4M/oNtuvY9rYEzX+UPez8oQa/2GcB8oWvzdIPfA8Xbv8A0SZHW8CUI/ydnfuZygQ8Z/vQ+zrtvCRhhF+WJQ0bwLM4+4xrr7sQYcMECYkOIitaGY4CTRtkMM/LZzaY1/Y1kE71ifwDnzrsQrGIksCHz+Tyjmtd3+xyBYKXU8He4bb2Lo01Ql8nYdCFtj+JHIsY5YxIZEJXoTbQmstuw6G3wiEWlk8sZ+L2F8WxjWJEMihol+I0bDQzld3NEssvuMe/0LWv9DHi0JdDdNDyPgNksc8E3W6y7new227+B+78DdRISMDtdiLcuw9S8jtknCHgLLNDbYxCX5Qyd/lDd1PBW3kgxNiMW1dAUVeEjIsKGQI1L/0ZsI0jfuDUNIWO1EmxCkpdcA7UWEPQ6pX8wlrDXyJrGV8slo1+CYGk4B9VlCaYEuW/Yc1jGTygiaZH7jxx+RGOY9zxEL+QVpbKY9C92+4/I0WqhLqIZPt8Mw+3wx99BPcdxnPrXkTkeBpfyiRBiV2/Yv8AsGmV+jwAVehj7tfsKc4oemhChQaGhlQhMb9hNMr9C+DTXJwCu/cd1MDRL8DYEJ0yngcsOZyd/gwEPtiHsSHTk+w63QTpDGsKQjd+w0yxjmpvkPQyyNq+hro0ayjyEUuW/wBi5QGvBFbyxJsQSESY5GXrPcXLkxBkWtlE8bwQSEiHYVtbKS5/6ZbSJNRlbf7F/wBgZtWQhBjbWUNX+cNbW5YuYNuf2PFc+Rr40JCQl0Vp1bGNUqNkKDy9IpKKDfx+RfBR1qxLo8iZu45TpUNwYHgpkP2/B7PwJq0ISEMTNDp4LuNfJklGoHLKSl/A/Z+DueOxaIaE7eQxNGsCbdOjHMj/AAmNptv4SFRKv4Q9GbfwhC5hjU8MsI0zPRjyO5SfLc9iitf4FSjbGOCNByJOJ52ETpBrZYYqatfyJHy/kqj/ACPBSpXCc3WxdIM9hfce4lyf5FyPyJ5lfkWpmuCZsXB4fWDQ1qYkzj7jT/ycDR7z/wDAz9fBI51nRjW7REemNpolTZFjNMnGRog0TpByGoanYN2FkbytjTOjD0NE6NEHMpmsf1qJCCEhrQhlbxDdlKjBsCELwleTIQSMDDfYatPLwVU1syibH4rRsgl0bNnBcJhj2iYL+B2TVvwOt4EqJEG4NilhwWWBq3MciJSIjyB6U3+OghLpBvsKh4Q3sloWOjlqhMqmBvz+UWzc4u41GxIQyPVhZKDDwahMyWiC5CNpb93Rm23n8hZEhnKF/aDboxE2/wC4IpFPkS7F8irKL5ombIlJrXVljQrGEn5yRmS+7Y7L+zFwkEJyy2+hd6H0YtMzHcY7fkp2ORSFh5HukxHAs9ujGhNrIojl9iV/whCm+X2HNR7R3A5RCCJ7fSCbeoTi0fsS1U/wXQ/wNkL74Fxn7INYJ0hCDHuw7TnIz4GpOJt+w1OSCd31g0Qgm8kymOngpVtshhYIeQ09BtY6MwL8r/YkJEGzUjb6I0oaUrNEJZWDmshCEg0RwMaNIs6HWNMd3jho3RtkJISIaKLSrI2ogVq7Ul0/kz2fySVH8jmp0QS6PA3Rr3r3ONhIYabWxEi/JfH5GrpfkyPA1x3EuGTo2JlJyKX+AYweDlBNErG/D5JaiTfcWg0Q6DF0Y92KxYUK0E1Zw+UXyad/MdJtvD7wt8ItwaNcRkPA9ofb/wB+x3IeDDeWkLCKT75HKR8CQWHwTiM+Cq/PB57HhDRPI1BlFvt/smo/CiFF78FUDJjP8C9MqhPlCH3MC614OOjwdoIYtTsXlr7CZLn4Kff4McG1bSytoRdcGJuj6NDKG+zt7mezSvyZYgOld0Z5efI/HfWGBipfjXf/AAZ9cGLanuOTT+SsVp96QWnX37dD/npOr37LuU6UvyJZO+5zKvuZ1fyYDT7H6p7CGs7H1YmaBC3zy/6OGoxrKXuJKYiGiGzi1p9zBGifK/2Q0NVoawSR4/JktFEijiwHrlvuOch1uQwQsiQlTQ+wZsSIEvP6E5vf9wkXX5NRYU80bTbuUnGQZRQxWoLTEIWYvkaXZfIgrS+RzUs8MQlw9HgbNw0p3JajSScoUyxpaQ7ZqDa8DaCoKZ7C3UJ88fsawMbSLbtXsxGubZt8r5HTdGPsPgi0+BVaml2Rz2EKS3r9Do7M0POBrFeF4JUQ0SAjkH4Gvf4DKUmd/A7Emz4g96hKfMi9xtKqbcnmYX40Os2jnEPYqJ/ANSl+xDf6AjW8/cQvxv8AsVvGWkza6LTi/Y1qOaJv7Dbrw7jGaUwZSabvcV10YvgefBFnbj7DHI105WEYCSwtFjScCiRvzBmV/IJdz5EkzXyPvEa2JrvOUJwsPI1HH03gizef0G23Xsc1RdD5F5fkX+rGpoe5EWT68HAy9zkaGiL4NDvMDQ2jyKI/IVg0+TEqnuSaGcGWhBlPhEGhBKIaH4UJY+QUHLxTv5+xTcQ1v0Jp6IJn5BknJy//ABEOjXYgpBmlhisZ0I5jpEnuv9jSCwVoZ3Bne+iE1fyXxijYiCrVCTNbFBET5CTuzRW0XyXDSHPjAkQYSFvR7GzJGcLBSWWBW0KvBRIxj19IPaoROP8AQ2YJuCS2p+wsWFdDvaDTs+B+L4EMcP7DHrEJMoSYYfsUsMXBvAruqXgUv5BeRz7D/wBEPyfBLCf4OayzZBa7BvrRGTuOwmva2Mki2Mx0m19j/jF3/wCQ3BVPZDGkq+4hu0bHOT5X9DeTX4GKU+NDnNnIGnFGGnou3S+Bd0VcUP79FfFsaxmIWmhfsdJ006h9lE/Iy7H4Yx/3Cfv+Rjk2Bz1CVNX6Emj3HNEWXAhqDMVoxWqm/cX+rE//AGZqP8y6WCO/5RWOL3Fl4PHP6Dzl9chsZIRfkrs+T2fkwQp7jYlfT7FEJJe5cCST4UMahJ0hlBDUg1aj+Qd9VPuYzsawS8G/wjTIl0Tq56hzGgbt08lEJsY9WiDoSZ3DL859E6tCbeo4AitPqfJ5RDcVf7Ezyx7QXTKiDFZBnt0gkQaG2nG0JWpZK5fQ96XkS8FRGKSHvWJUSIRED2Dv2Fqlo9sk14JZrlH5IylTHWfWELaoqmd12FJaRr2ySbwhUlBPY9j4H4/gQuPwPeMQl1LndwxRNl+BR8jIgSLD/B5fwPzfAmZs17GHTqXWCa2VYZts7P8AJD2bfgZCRCU/AQX/AIEhPuDKB4dh7FX9+hMmQ2HbzXKCJdZwOasMzETFhad0cEn2Gcdr5BHBS08PsKa+Ae+sCwxjVFNJp3sxeK+eLkhh/ILz/I2Ym/yPaF8eVyUcievBj2F+RaJ0YykZQ96/ITf9Cf8A7HT39ymbQuTyY1UkN/gSmxjIQRRqoalSfIm7Pkb9nyPbjDWlTTEq1/Ioz2J0anVqqE4pKW+IopCT2ZwJBjSxTok6wnSGAttZwlgMiYtjd8CaYyE6wc1HiJt8v9jSCxttDdkH64RCCQkQ0NFRM4QjgIaCnAituI1lDzz0QujiGGm0QpEQkSZ4g47FphjKPqunuNNtItjtyw/mm99NXcofaD7AtkqEhIS6kP1ozWx2MHkVWjY0f4j/AOM0ll7GQ7LKKxLo3gaeCEj4CIGIk7cDVy/gXxXwTGmaGHRX2EPa37iQ2ghsdshLN9S4bY3INj2Vxp/ASu4U9T7hCInsRM2JBiyqMZKtfsSnEncusE0k3caETQsiJO0JbWgXI11ergOJxVE2/wDIVDCyJgO5DPhY5u4ZCdU4NQk9r8hP+g7Syp0oMLYYlScnI0NDXVNrQpxkpm0X3G0cKkkvuNJmnsf2iXKGujXSdYCCYMZ4k7lqpMcM9WyvXVgfRpMgduTlmGqxCxY63WJCEhLpKJWJkzughIVuSEb/AGJaGQSgiCQkSDd0OcBZzQrmxNFv7lrEhaZQ5KjmpOs6N9yBybOYLENco+ZobgGwUcP2NsXRDGmpeSa3HJXgj8A8NBvaMQYdo14GNpXgSF0eIVQ29FUeWYQ8ZRLsNEL/AALPH4k7Z5g3v9S7WiGbCRJORoH0SjM0KvgaJ7fAlnkif9Q+Rn0S5INJtik2hjcDQnB1r2K1l7jSfZdGNA0M2I8HwQq7mQbWh5CZBjEMbfAnmKioLWw2lyHw4jypCqqOBqPOydIQgwxb+5tJx8bESxuI4Tv7mVAipGo4xoZOkILwaWtzN5+Ygmpv3EMJBpvYJtofWdITsJzAiif3MIj7jdcggNnq0JrQeDZCdFLJu1j2sQgkJCQsSsFtIQeSRYRsAWZkSqmPa2QSEidGeTE4uYnWHKCm8SSJxpd4/oVESAuiRro2uRKMoQwcbG7N9Cg2LzEkYxp6EhInSTI8INPuPF0Dl3GpqzzQ7JQBjFSKyPPIhIaSQ8ibQzOPIkSLq9LZkRV+hWRh+DLC6PGjfcSbTFHExm9bGqzZrQ2pGx+RJTAlHxbKZp0I4fwDt/5GiF5P+IJmSfBLTvQ4mt/hiyYIzJ5W9DyBK4h0L3eTBpX2HaRPmC70+Bd/qf6UWaLYoPuLsxOklWyjU0LuGJkAtXHyU6go2txd8eUZgsccMLkeTBrfldy2t6TpOiY9K/L7D7TF7dKRTCe2BFOSDHqVX5vkWVSdJ1xHHI2UsmiYqoFHchON4cJNyjnM3pjsrJsaIQglXB9PPP8AQ9C2xs/KMkqCRoQ1WCb3QetqxXZjop9+c+TwyCQl0Y8IJ2b4HHM2I0QmzlhZUWoceeBM1WuRCzoxIguiVsk2hFi0ZL1SmpyHM8sUZaOat0fsTQlMEIPA/BDPgiEBGuT3M+4b8hp2FNvKeRb7j8DaBdG5scrFRg0iXcbp0jFKuyLzGuTkSlWp+WJWIHQCV22JwbY84FTeE0JNoWTRfc8iVW3Y1CqHyT9xjU/cJWShjaRiaPD8oSnTdY+4tDNDtv8AooLMbVqPjUpKW+3Yxgq6CGUi3gex8GLUU2ToeDIdtf2PibEORRRZewmrAQ/xdA40jMQOHlPRUxDGXFOB/QjAdax3TIu5e4J9wT7ws8lD7UNRim78MbK0fV7RffwVJYJo1kyBFC8FF2Y24aldYg2w5PuTD2E6qusEm3NhaX933YkjKOUWA3cRZHgIjafDsytVr8obY8Caeuk6We9rwJmkTMeyErkvNqJ8BCWxCe9+Lp002PXQvzv9jlE7kg9goYtaE52NF9Y7qBHaDt0hhWQaEJ8BKjIVaNkTopbNjKoTWYROx9hsYM3rINPaHFna30wNtFAPXyf4RKpJl3al7Je2NPA7iG6NYGXMcf0NNo9l7jQrm3wO159gv1Hz0n3mDmhl33o/mI0VvYEeD6SU8Qm2M6cnL8DRqJHdB92N3hnZGVS19hNgZPBib5AVfNe4xyI+i5P2/sdeWRtv7DoDdA49bn5EwZXAsdBKNpDZm1r+hcZGTjnoU7rQyzpwLvgZ7c8mLzN+BPiSOSScykcmhfxB/dIPUQ8CS6F+WNuSZgMp4GkkHdSLzEn5k1o2AkYT5vBaNdmNjlIJNotjpfmZFro91GOUxAkw4ZCypE0x/ormjG+jHwtvwiGuqeZCMUlL8ThqP1H2OzI7AG0E6YEXF8LuNtYLrI6hjJkEcgdJRAlQbRGsMgW++/2Vw1gaS/cjgKnWPIg+RTfgVWhdx0oeXWJdINFPxCbWGaA7IRwGaJjYo9wfkETSTo3csRCCbeoUktDG1yMWBcLlqVGTdMQcQcKiOPQaayJqi035G+429iRKNo7IaxXsMyux+Ia7Ii6QwlTMBoIaLoV8G/8AwVpxlYhR4ojgV+xjNskazvca7Y1/xDVf1DCJKfEGqb/UNKm3+A26I4bD2VY09CMgXm9NmUYzZSXuZO/oKPH4jsV78C/4A1gn2hGkNWYOoxb7/wBl1o8CaQbsC/2jU6IN/dBJ4A70l5E+2J9opwM1GpSqjVuwd2ycBqgdOal+RIbMGgeqOJmghFYTYVOi7ttKD/cJaAbmxv8A3ojMfSUY9YqGJi85X5jCllM2dJtszEwbyMoXshV2xCdGqKrKYijkz3RtW4q6qOxzGu0yuhVwEWeFoSJ1hkWbQWzJkbovLtEnAsX5X+yORGEEGNwnrY7kxFkiybRg+CdEJUg1RBu1OTmY5q9DurGIrAewN9gwOQxqxCEiCime0KM5FJsSJaGbbZjLDYgqXtOiINUbGhj0CufAvV0yxmpmHsxoEh9wPyDc7FEoXkQzIhDJ9EF1uP5XcwJuRbcCGKNYfk6I+oKPTDtgktu6IRKMl7un2YkUHzDc8L9mhk7DfsNpyGdsJOU0FxsJq9jgMcE0hj2YnjqERTL2SD2MZEiobvGldLsJum/Iu8/In3PyJ9wslhipBSjyQuFb/BCRDRp1ENEFUVkhNXFswE0dnWVmYQi6HVGqNXX04HVzC5Gxi6SkQxKhmGlE+yJuUcFAUvMQhwdt+AhPTlaEpCI/Eb+JZSQW5EKhaRjTx4EqQg11cORI/wBCE3INJI+hhV3f7GPLMByiJokjWCwwi7se5J0gkQQ3GZYhK2QYqSQmJHiF82Hl9ITo3DuF8hjp6LQmvIqaaY066NoW1VZwZCXpCxC8CRBxTl5HpdldeWIWg0y0+z4Gn2fA1BRfYVzjY8BLo0NpWlDhWOZjFoqRcSeKjdgbbMjTKfYptPwKxDohEq8F2W0a9IqeBjZjwp8ofB+SEcT9DlP5IXN8iE+0LYyYn2ErVYFTn7CmivaGmh9H4FBpPkbZZW/sSxIl5YpZX5PA+RPt/JA1XfIjY8DtzNCchQ1MGHSgcaM+M+QCbUibtECjtGxdZli2DmdGTuLGBkING5CClNdlUDmDozt4O0mURT5icYJer6Tpck+BFecaiGNvBmaIg0nsfkE0xkGuiINDFcBJU+guvl/sQSSVYjwwO0kGpaHOoG21foSJ0b2K2iFBrTkjCHhBnYftOAUbbVi6Q0MNgowxzR6HLnBFRBTUTyNXqTtj8BziTokRJCVO5Ca4JHeaDaWjBNJYYx9oysD3/wBjltQwipCQwk+hxlFCnliZOWK6Dy4PnDXMdD4nY6p+wLuBEjJ1iQmMkeDPt4bFrMaaHgV02xexUmuYJimc56JFBXpswmu+SmJCgnB7Q1wNDo2I1XRUatLucQtWRLtYl2sW8JizyF4h2wWF0Ma7EVGPCkQZE7kbE+8XvD1hiCgRVrgq0wYd5FcoaEmmYehoY1yVSVC3h54KEsByrFrsiY2sMZk0RPKM6FljRCEIX110A9Us08FzVAnw9my+R2shBohkgw7kPhQvzv8AZjYSZwEqwpGklZxqeBIQ+sGIlE2C9BuKLYx3RPpLHjLG8v0XhDXRuKM1TRi49HfBPFk48jpyPkppDvXWxZyhK7E+GO1qICdCNttii2nRdwKMsJ8jupXHplmqkTdDdOCTeWLBofgVIIO0px0wMtNJ9KNjF3KjcCC/1scISQhDZKpXwNtBqMYgYMMn4Hoj4EmC/Yux+DNUvwf8UclFdzUQoOUYT2PIxjRHWbHoHwQwDFtS/Au3+BVyg/JRwYPwxHpwIjLCH4GhoaQ1UE3AMkSupKCfajupDfgV7EMKGsjQjPIPcGG3oJ1dYLwd8uDfGD80K6w0YV1PsODtx6E1wJRmnkZCDGbDCIB9oOOpR1hvuKKcdFhVj0bGiEIQnQ2juxk1rMuGI8BzVk6TrUtlEJDmrEo4wOq2sboeZgkRd+iEUhow0Npk5QkajoTRY6G+AcD8DbJ8DaNQgkbwJQhe4uc0XjTSwID1OpT7UT0vwV2nwI2WUSEcqLORdNFriGbJpuzgSaZ2JISUH2tDXchw/wDhF28GRyT7CX/RCSZsSacEhOGF3GI85GMTQGO8i4O6vyM6T5FRqCknPycTX5PE+SzBr3KUni6NYE4bFbaHF0YxieYqLUrmPlmTGBRUq+5Hj8nKOvROq5ditD4pnqJi1A1BjE46PSbYqVNSIaqEVJ2MnS10K5vNm+EdznryS5HBG1R9KaCk8BI31BrOldiYm4PRkMucEydYQSdiFkjx2O+x3AaHsK0XRCDZSQbamYHE0SkIQdDyPgaVQY/AhUnPTZCEGSViVhRwGWxLFaVFigsiC5wq8DRwIs8F8pbIQg+qn19x516L5JYtGPMP8iRvqAfAOy/JdmoQj7nuaDUIIajpRDjETtbwhN3iPRP9jH2HyMf5nHT5ITf2Y8BLFqOs5Hmu+RIQzKURyHgWPkpLbyxRXR9x9OzE27CdX3BOLtkXK+jEk537/wCRMQ17nYRDI3jkZcEn+RUUGuw+++DvMIq9uiclWp5I+6GadsdLpkKl5379EReIi4GMzeeCOFMKzN5HrryJXm4h9xnkYmumx+4YzmPjVsjW3+xlOfI0PoxjW9l7j1mgQWNOpPkLuDzhd0Pu3K8VMo2soctbQ0UaDz0e/PgRrPI7Kq6XsZHSZ5Q3yBNNMTLlsIuxCosGlakpCEIv3x/ZyMxlimi34GgCc9CdyPIQPaEZAmgU0NIhCzOWN8sWA6yaY4c6IgvcbZFmBZehuXMSuWMaNBLQINFxstdSeBofIKarTIPHRIazU52NizFSbl+gtMdlgu5YgTIDZjD6ENsTVmJ9oDBuIeUeaN23IMuPuR0ZgdbeB5Ew0ex9gip4Y08QlGhmNpfsh8EZQDfOnujbdx1uicaxPkmeYZz0Fu0Bu7YQ6Sb0TowIq28L+xtJGyb/ALE3/Yi/uR0GIoqP3H/3DVv8xCtkop56f7GzNhEp8DJoUQx6CrtFhCaQ2h7mo1upBmsKfA+2OP0BdF1I4BXqz0U0mNPo0J0cwpfbEQTlVps7EzWPxP8AQhf8Iv8AjP8AShv4b9h5Mog/uAyWjU104CNCcnGhYQg0haGlPFO0V2m2Z+BTFH2JFwxz+5Cl2GK4sT6PBiuOTLLSwhMDRj9BZVoyNf4EW2wqwO8QtacPZRmmN9ozwTpWfu/30WCyHzdoT6RwtizrIqGk1wVMGTRuLoCTyeUaXYU0166CJz74NYZs9xwQUO0E2diGUmfeXzL2sfaZHg6LAwNZtf7ESdJyhVuahUTP/A1M8dYmJnTWSulVmlLITBtP8HTDE61AJrWyNqRmQ6JrPZBp4DwCqiDV7j7AXYfA8mGqJ5udvYWRzIwzUm8BOLXAsI1kR/xF/wA4iv6jK0L2EKhewv8AnO1+I1/iPuB7GeA3krZ4IkMMXvsPsJRYGuBBVZLwP/lHDHBNZSXgXH+In/4n+1H+5CI0lGO4znkwGNQei/DPYgiGWqHYSQ/AeAT7DwfovYIjSoeX2JCMQY8ZHef+lEC2GNDOQE4H+9Fv8CwjwHyykPr3IcxN54LKM3jKKSjNXJ5f9C4EsdGhPV4J/wD1H/1DK/uZq2vkynyC1YewCTYgpt4ySvvv9jU6SocCC4tDG7wIEoruBKwdpRJ9I9h4Rq4EPhjol0bFh1Cwl09lOHYi8irPbGqKpDWfR9My0Zgb1J0e46GpQVjUxeRtIKpNcclja9ew1bIadvTalxwM8n4GqeBBj0DokJl8Qqq1M2XLB8jq1l6KbgmSX4n+hDV/iJa/Ef8AyHBX2Gka+D/SiB4F7C0QeZWDT0OqnIxFd9t7DGjGR8CZ4GNvDGd0jhMS4PExq4YmLTM1GhY2ntFudMeWJ4RNQvtaWurboMao842BajJ5vyLkf5F3PyeX8nNfybh0dL7Eoq8Ie8Zm2uSxw0vbqxrD2YaycfkL/pP9jMn9xf8AaNL+5Q2TJ3CwNinPuGU3/wBQkUaBwNqwouRAg8w7piQkZRCfRJGDGm0eiUfiPLG2tzGgn0g0RtUI2mJT4DHEccDAN2CUJyZxCKdJV99/sdCDbkMJUdZNMiiGaYtzFwKJpRGZpVFOFEeBI0bZCC242LT5kVWZh6LKDMn11fQH/wAg5ysE4JBEwNFrqevctY2KSUJJtpbg1CD/AHI/3If/ACDR/gQ4/AeFQvgziZG4SXokcDQ6R82vcd4ViPwfgbMaWiUa0NnA+yPtj4UPuPggNWh8KZThiU6MWELI0LbYsr+hZtop2gzc3I0MI2H3vyef8j4n+SnWPcodfcfd/J5fyLu/k5P5FHaLKHNm/wBCl9wJOj/wEnVkSo2Pi/My/wBzPqbFtn5PD+Twfk/0MX/QJHH5OJT2d5/0Ko7SqvJ7EhOrMLTCqpB4XyeELshK4DdwEOGBb25HeEWXcLNd7YsSdIMTSYGhLZQTQ8e55fyU/wAj/cxjP7F1iafkTQYRiMGQksmhobyukGhrNLo8KBi0w+iiuhG8YoUy99jwqPLpCRRiJFXOjVpSidwIDUNFsMfWCCRoYSINDxD2wvghKFZJjovCeP8AB4PwP/mLTCUUGiyPLr6INUWZForJljn3tsRaMHiH2B9gfZZwUx38hhEwMMuiXSCbDxED1gwQrHsgabRwKPyD8ojbLGn+T/SkJu/PoTbWw8etNDETDQ2lgozeBs/yGv8AJjbx+SDDPcX2S9yv+R/tZ4/yf7WJaetiUX45EdGxWx9jL46MyKSrkbuPyOVLGJCoXOhXKF9nSSh0E69oxZe5nDXAoz6GQ0MsGhbUWuZJ7fQAGwSrsEw8Cq04N/Mg4GMryNmUJrIuBhNV+R/qY/8AoO/+R4oPAkG+SZENCNvAo1V0YielvQww9R8CU6YjWTpCRaKfkM16bL0GgWjdC2IZqha66C0IWxm4tdFnbouiOeqa+gtGp+EfuOWLqh9Y+TZ0Wuuw/QcOvMeuiFs2D2PpGPXTZn4B+IaMWjQLQx9XTotCNRwcM/IN3R7H00GnQPofTkZ+k29YYzgYzg19HgRyM3RobjZ0+RjGPRoamrNJsPY9mk56OnoZj6EaCGbGounjp6dP/8QAKxEAAwACAgIBBAMAAgMBAQAAAAERITEQQVFhIDBxgZFAobHw8cHR4VBg/9oACAECAQE/EHUwLxnpHrC8Q9Q9Q9QXgHoHqHoHoHoHoD8Q9YXiHqHqHoHoHoHoHoHoHoHoHoHoHoHpfo9A9AXhfo9Y9L9Hpfo9Y9L9Hpfo9L9Hpfo9L9C8b9Hrfo9b9Hrfo9b9Hrfo9Y9b9Hrfo9L9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9C8b9Hqfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9f9Hr/oXhfo9H9Ho/ofhfo9X9Hq/o9X9Hqfo9b9GHT9Hqfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9b9Hrfo9T9Hqfo9b9Hqfo9b9Hrfo9b9Hpfo9L9Hpfo9Y9b9HrHrfo9b9Hrfo9b9Hrfo9b9Hpfo9b9Hpfo9L9Hpfo9L9Hrfo9b9Hrfo9b9HrHrHrHrHrD8I9A9A9A9A9A9I9AfgHoHoHoHqHoHoHqHqHqD8Y9Y9KPWafgvgvm+F/CpSl+hfoUpSl4pf5CL/AArwn/AQ/wCPS/SfMNIuV9N/FfQpfp0v0KUpf41+FKdcp/ytG/qv6DKIvN/gv56RfBfKl5fF+FKUvzv1aX6K+nS/XvK4ZfivguKP+JSj+hgo/wCO/g+dPxX0aPhfQv0aX4r6NKUvxpRfSv8AEpSlKUv1aX5wfD4o8/HJPnfnfqP56f4KcKX+PSi+jRfNfSv1s/xr8m+b/KX0H8H89PC+N+bKMf1qX+Cviv8A9i8X+ZS/Qvxnxhg08r5L4UvDYlX8r9KlKUv0V9BF+S//AIB/x78n89PNL8r8cjNvo0pS/RvFL8qU38r/AA5/D1xRfUv82j+g/k+H89H8Bi2X6i+jeV818bwn8l9Sl4vF4X1X9R/zZ9N/PXzhp/gMS4X1LxfpL5p/JfyKLhfJfwH9efVpS/Sf0H84afjfotwo38VL9S8X69+K+kvhS/UXwQxF+V+T5f8AGnFKUv0bxS8X5v500/Lri/BDxwTGJ/K8dcUv0r81818KXm/QRfnfmvjS/Vf0Lxfhji/Rb+vf4ev6NLxR5GhoYwvp3+ReL87/AAL8qX+A/oz69+q/i/pz5Q0fVfxE/rX6N+VL9C//AJVKUo/4tL/Nn0NX14NCwLfLE/pr+TS/C/w79Ol/gP6dL9d/wKb+erml4vzfDYxQ1+VKXi/FfWv1b8V8qUv1LxfhS/wX9F/wdF/kVmr6CL8Wx8Nfwd+tS/URfjfnf/wdmvpP6l4f8O/S1fUvxeGN9NfKl/h35Qn10/5r+k/pUpS/xX9LJq+s+XkWxMv0ehfQRfpJ/wAucL6dLxSlLxv4Xhv6j+gmP+VfoPnV9dsbNkX6lKb+hSl+ivivnfrL53ilKX4zil/gMv0GL69L9F/UiNXN+q9FE4L4U39BOFL9FMvzvxXzXD4vwpSl+d/n0f0H9WlKUf8ADvw1c350T+LJ9Ey/OiL9LPzXyv0r81/PYn9V/DJeKX5v53h/Xhq+d+N+LGN9KlL9el+VL/LvNFzSl/iP+Z1w+L9R/PV9e8NDQsCf00X536K4v8KlLxfpt/F80vwv0n/Dv/4mr+HaJi+pfoXi/wA9b/irii5bKX6dKX+fR/V1fG/G/QfCLxSlL/CpsXyX0F/AT/j36lL82xMo/wCLSl+teNBfjfjfm0PBSi18aX6N+jfmvo5KXm8X6N5XLF8l/Bv1V/Fv8DrnVzfrv4FoT+si8Jl+hflf4S+i/heKUvNL878b9N/xKX+BSl+Or+Ex8d8IJ/Oi+nS/Kl+VKX69/jUvxv1r/AvF/hv5w0C+tS8vhjb5L81/MX1UmxO6POXK2QViXcHQQthCe1BrYmNWmNXQ1bX85fTvwo/4GuGUf0tHFKX+BBoaGiwsX6F+muF9e83mmkMdCbsdhiXpEOEaViVDyxElCQbCw6OHUNVUWEYnHGNNZ6GuSR4nCbTIaRr6I1v6lKN/wm/4PfL5bF9Vo+VL9WE4aGvgpfmil/g0pfhGxjSEzoXcxK2OihdYhekRLZGHFhCjLMtgwUCR1jyNRJC54eUhODUZI9ic2NTKMPZlYZPIw9kaIhbQbtDTpj62NXQ9xfG/Ol+k/m/o0peKUo/qUpeKaPnfjfpsYhOr69L9Dv4xsWkhvoZ2xJ2xK0hdQ+w/ZvREnWRsi0KeSzCFhWN3QoVY22xKfZDBIJG4oajMqiCwnZrRIqGg02hNPDGu0VPZIYeyNGGZWyJ6Y6iUa9Bv0jpsb9MaRPaGmt/S0UfN+vf4d+ej6F5YvpPhBaEnxv1aL4JUWkjohOthLunRCWhEbeDCIw4jIwjIiWzLIttmRGTHWJMmU3kSLIdashkNVFVo23kVsN18CDBoSMVTp2LsWMoeECbRlkKoaWmxURehkQIxEyllGHtCT6N7QvAx2heQd7IthvYbND8Aho2yGy2uL/Fb/gbKUv0ME+tfhfgxjpRr9C/RSbNAhM2oJgR26aALSSR6EfeDAVZhbYm2H7ZHSI3sqWjJwhtsx2PohOzDCEmzHux5YoQM2pQNcLRBqQRmNfGyNwhqoyGJiMaENaE2soizRGVYMbIXRjJNoiehpjD2VtFET0ytbMMjWirtE8M+wx5MlJRsH1oPYw+hifQ9pE+TKUReLy/5mjhO/wAG8NnQ8jY39PeNCE7oYCVt00gWgki+jIiXYvSI+2YWjLREtss0RvLKkVvCMdshaIEWzo2eBeZhgKtkWQYxMG9FwhA1USokxELBq+NfHZp8NPA1VBBumUCw8EX3lITmGNdhYKthshNrBE9DTGWzPRWsGHspZR7ETMDHZPDG2tmGR9DflGPJlFS2Xwxq9pMbth6Tg1bDTrPCG62uaXml+V+k/q6OaUv8JuDd4eDJl5hpkdINBHbvCFopF9DrZh2XwiNtmEJvpEfYwitow2zDXBEthzoQIltj8BMJ7B0JnkxoOvbGPZCxwXZjrC1wkSB7GQSa2bINYfJOFiSJwnB6TFjaXDzD0NQQokYxoq22OBY0RabHAm0RoSC8iNoahfJD0Ro9iHp8FT2j04K20ejKmyp7PRjbWzD2TwxtraHRPDKmyBx+xsGtYGAR2p0g9pE5vDYuaX4Uv0bxS8U0fKlKX6zYymbIOkh2gjsJXVEiL1GvLKl0ZekezMLSK2kexhpGWj3FS0it6PNmGkVtHuNGsjZ6E7yeDI2YnejHsNmJNvBFtljb2Ez0RbjHvhIlDGzwoBjXizrGMQox214SrnwEyQSM0nz+xENCiDwfcqeGNNOFKmIZ64TTwGnXHgyJ6GoexG0NNCYyG3QmWCttFdCbRU9oh6ZQqe0Q9MjFXZloj2jbKHCPpla2ipkumIM9oe0hkMabQ2DRI2QaNr5X5sXE5pR86Pp0vzSb0LQR0gx0CTsLzAtYRhxraPYYFfSKeyILwRQhsTS0jLojsw0imJ2RPY20hM+iJsb9KDTbPxFWgbb2J3knsGz2KsIkHWFjhrzpELAgmeEjH3jd2YEQGbcJmNy/s5ShuvnrxRqy4pBjUeOEzGhgqE1pjUKvIo2NXI+4nNMqY1CngyHpj+4m/JkNNCZdkPZlsRoTrDMBsuxMipnozKPYjFLRWisQ9MwKntETKWiuzB6MwL5RgyP0HuBu9cIS07wBp2h/G8ofzyaPqpMWgOkF2BbwaahFBb0jIaXZUujLS4ogvBCBK2YXRW9IT9iSey+ERvoXmY0RWE76IbKWEiNhTshaQwJn0QhhhCPtCd9E6KNsR+BY3AcaEYmeEiPcMe+NAhuIMmTsDPlpFsyyCVjZ4yYpsnCNUycYMaacIQyUJwhiXCJxrswyThNjR6HT7Mtwx9k+E2uzD2N/JnyJkRPTGxWuxO7IfZGhR2OM9WSbKRj1ZkQ9kY80VoqfRG0ykV9lboh6ZEL54Q9MbITEPY9hIYDZpnYHSG0Q01v6ej5pnpGkHTHQBEOkotJENF2J8lPQ2ZbEl5KhW0X2yJtkLRl9kdsxI6FR7sqDvQmZC2xI0hsxM9HcZDSG7sV6Gt2zwWDD2IJuLeioaz8gxkRU6CG7swVyyVhD8Dgl5ehLwlgwY8CTbHW0Y8GPApsbvRjwY8CwrB/YS9E9GjjwfgX2MkwR+CehfY6OGfBPQsPQ0T0fjmPwZ8C+xnwR+DPgz2hrwZ8GfBbhofgZKxO7Gwj8CbWip6DfojQm1oqexv0RrZUQs7G3TImyip7KemRC9jDG3TIhexU9jrTIFFTMtMgV9sy2R0yGitbKhpeTwMrWyC3sz0NmhskMaY/EI6ybIPcXx0QmekaAbxThGwU0YWgPSexg9EV9I8hER0it0NwhbLNIpgTNohbMNIYJnRhsYaQ2iZsx2yzSG2Em+i+ypaQ22xJibsjQNmzOhdmDoZGwbYwflY22zIjaMb5Yz2ZkjYtjGzsz5MiWwbsI/JGJNbHWRrsryJMZnyT2Z8jGfJfIz5NEieyez8j9z8n5PyLUPyfk/In9TXE4/I4yQwX2VPZhlGCpFTGWjRSXhkbTGksmCFsjHoRIUGWyXpjUFBTaKaHAoJe0ZEdDwe5W6IeiNdF+Cm0RiuitDR7XD0K0e6KFOjAbIh7RtA+lB8YkJNpf4JakiyhGMNswK6M+y+2Q7MLRl2U2yG2YaK/I3dinYnmV0yN9ieZZ5GXwO7MTslbZ6DbfZl2V24JKN+yLyJmTcx4xYHH2KtCRZYhB52yLzwF99j7GRCrXENWosEXkaRXJCQYe2RCSeiLYbTyREQkQ2njhgSRgwRECSHGQQJKkUiXDBjkYFBpFXBcIjHgiGvBh8Y8GDBjwY8GOMFRUUw1gbnR9gp0hI98Uplsieh42iiCbbR6H4E5o1yjLQ6uilFT64MropGe0ZawNtmUeRFT2iJ6Gk6KhXaMP0NujDgy2iHwVTyIw+iumNKyrsr7XFPRF4e/6X+ENsx0ehHsQtsi9l6IrfZmS2zEjo33xjtkNIY+yrwQtsxPQifYrJbZU0hu7YkheRF9j6rBjsST0bDOoh9xgXQR2ydJDBgRrsZOwYFHoS7ErCDa7MCSZ2dj7jBgSTKhUzHgq8CSG1ox4MeDDLCoqMeBFPwY8FXgUG4Y8GPB+BaMeDHgvoo/ZfRUVFE8FKUeMotKUpYUpeLC8XjXFKbJDJSs2OorKxN2S6HBkTGW0TwOCsgW7K6Y4KEGGNumNIXoX2iJniGgmhT2iJjKIVC+UNGPqInDbtGR4iLw1+2v8I7Ykp4huislbYkWnQ49sXgT2zHPBpPhHbHGkNvsVCojshpDfYgV9EXZPSKjDErL7hu8ChjwUy0fkHfCrwVzMF1KjvZV4MeCuWscA0byY8GPAke0Q0VeCrwYItsqMGDBjmlXgb6RYVeCrwVeB5L6L6L6L64bKUotF9clPZSlKJx0pSlaP6lKWFuDOmi+CjY3cMrTBRRRaUrKylLR1FKE2WjqKzIm0VPY2WjJkSCp9DboyZEgw9ovoaQyIKntGWmMMiQVPLRHTGgyhIG/KIfY1EQSC+UQx9REExWPc/S/wzIW2JKNFot2xD3ZFJWip7ZFwi90haDR7ZgzHO2JCwHsbMCrRDbIaQ0e2QJHoewJaD7DAknoSbwElEH3GOCpVibsD7uH2cB9Qjbh9gknpDWQavZfAowYXQ2vBHgq8FXgwYRV4KvBUVIXllRUVGBOulRV4KvBV4Lkq8FXgjwfZw36KR4PsG7opfRHgXoOJBmlCmBWNibaMTKUptVoVFKYGnQrK+FG+yiii2NmWlZRXDwZkorKzLZvTHUUUJ1sbT7GkKWxeQnIe8EfTHBRZntET0xoKxNdlPZW7hfTGkKxdxD2RPTGGAlGW0VHV8L/DLbL64EjbMLSG27PuE7MdiJ7K+mU+yzsJ7ZZoab2x+4xohbZgG29s+4+48myr3Ru9Mi8kXkXQdgQsYDSeWyLyQ+xd2y+4PyYk8kCVncHWEyLyQQJdlXRF5IiISESHDBERDnRgS7EEESFGr0YIIiCEotsiIggnBDrMGDBjjBEYKIjwZgiIirwYOoqMeDHjgiINAqKioq8DVAmKoqMGBpMWgVFRV4KvBPBgwY8GPA0maPwfgq8FKuxzopV2N8KmRopRMhXsw9MaTkspsj2G33wTo+wrD6BtrZRIJe0ZaY0aylorsh9G9MjMq30v8MNZLWkNtsyJ3RC2KlpFCMSfQnE9ha0jL2RojZXeDDQ2EZQnEbBq0H2CTPQLQR2cjbhKFFeChr2VaB1sorwULuG0whRRRQlBpiiihstkZZZRQ1HBOiyyyx5SXosoooSmKKKKGoqJh8UeF4fdw+4+4aiez7j7ieyeyKlJ0RDSJ7IJQdk2iCH3E9kQdGLyR5J7GloryIU0ZCIggdRhkREREDUMGCIwOcYIjHDyRMgaRhCRaMtkdEdkRgQdbI6JDBUtE9lfeCehqbQ4YaPdGeyHoaS2jBgf+Nf4Jgluyp3THQbPssTPQuwqd0bdDcpiZ6FtbhD2N9IooTbErLwdTPCVlFY0rgdHJtBWVlbE+3ggGz2VlYqJtslYFb4yKiXkbNmeM/NufcSDJy0Y2Qe/hsaLAkkpy+NITri/OcaYNq/FKqhoqJxXw7LYWvsg6uMjW42VTsyZ4yPsti67D4yaJ2Ycs8TNNG9EIyMjI/HEZkjMkGyKIzJWQ+hyV4KZAmpE9obdDfwV4KEkw9oy0xv4KKE1N7RPAZL+F/g+hjae2ezEk9CXtwSZ5GvRh7ZBAkZ5GeAbNlNKAmxktBtPLfCBI9DQrCSwG7ZTRfEguAtINmy8hJMrBo9l8D7C+Aq6GktFRV4KvBjwY8DdwhNLojwQuiPBHgarCWREtlXgq8FXgq8DRKtCNsqvBV4KvBHgq8CfpI+w+wq8FXgq8D1pH2EeCClHrJCcSLwvC3A5Jt0UrkoqPTK+FKVjk+4TpUVCiijd7HXsKVlGxC5Lgeiiiihu4Yk0KYKKyspI6isrKyihMrMlfnjPni+R+DHUVlZQmWzyINumMrL7F7jot7CJsbfkoZozPQz0xulePyZ/aQmei/Q9VG/WCsvCcTcyVoNti8JnoU5aD0lGdsRONIdpRvrAeeUhfYI0jb24yRiZigbP4+Qpnmcb18YP8glM8QhOMepcJcwQt7MAQnP3Kn9nN5hLLGSYLxjV5eaextPXNXCKFFUbKKnplXklKtibpkeRTTrsTlYPYewe8xMVTE2Ccn8ifiDxM9w9xlZDWziyBll4iGlxvI5sdbyNG2JumQQJsHkbQksNkE9bjC7E5w8jcVEjHtCyEQNEqLUG+DVsqZRkhCH0NpDQ4VFXkcPI6WieQ0hKnsxOaYkeHkx4JJLpGK2Je8iZ0Jt9GLyz0CR9EWXk8yKaRkx2yRr0PjDyJEskvo6FHZHgTtTo8D5WEGJZdH6FPoeRcFccAwmjrZk6fYJ1TL8DVIbfRDEKdDFhbIuhY4VjutEJYjyJtDew2KrOsbC1rGYyJF9yjXkY2Dd4yzHHR2ISIrGg+NkCRk1U8se3F/orKxUWybLMFoyxGxyd3eiLhi6wuImTKOQuZ5pERGreH1xF4GqfoQjbJEKDq9BiSFQaeGMkq2iDSajE+W5SzTTE8C06B234j4eVGLeQjBlFkDdovJcHgykUPDKL3FoeUXsw9ncK4e+EZPZ5BejDwxKCfk0IeexZGmip4fBrZBMjIbdFJZEpD0NkJkX0DZaK7IaOgNWiRToy2OwJXodJjVlcTyPSMsxZ7jTSM6bbwQ0W0NG4w1Wg2CuyprI3YEwkWxotIbMTPZhaG29iTF6G0VsSbGkisZsG6kJdnrnLJwE2Q1g0dAQtcQx2MboJLBcZew/NILWkjELAjUW2b7LfCErGMfgShOLTDJ3M1kuKXGuv9I6Jxmn5cIxfR3cQwYyyGpcziHZEILREG37MWcriwQnwkNiNTe1/gpxwpjHtSINYyOLp/hJ5FELGN6DoqeuGt0p34BRPAjyWhLWMic1sR15E/JnhushDxgxLwPsEcNiFoQ1M9CzAXgJ2JD3ghlDdo9CU7Gi5nA26KayPUggrGHtjiEzyhBLCFyNO4W7Y1mBj0dgm5H0McQJemR+zF4Yn2fcaV0h7CGzLwM7GRNwkMErukKLSPcS6hdQl9DQq0S4wSM5ZWip9DSqzwDPQ3iV+jNH44VeCN0OjwJQ41xIeNivIsJclKn0NFgaZyE2kiL3MVrN9cqh5edCjSMgCKyIIWITY2UijRFDl3MhNs4owNl3cVi2MKvR9EBd8NCp9IWBZIm0a4el/vFGn3iJEinQl5AxIkilNIvCtrBIcZElkWlzZ/kJqe0MiYqey3nnILaJvYW5RfJBpGUKUnG1k8P4H+QiCSMd0PTM8IIzqAIKuHbvFJxDrQRz+S1VMRbImgvCGFQxrjwJbQzJRgSjPGSkfoa3YG1D8uFNPhrAlM9eDwFx5E0mQsFmjZkvk2aHtqvZlaQWuJH4CjynxTPLH2Gn2R+holPUWp9IbMKR+QkWWKczjXjoSzkb9hKzOMsbWTY9aGWsTViVlbMeBDEnGzDt5OkwMYmIgi7HyhCwjLLGSUJY1gK8OW4NnoQRhtnQjwJJIuNDcdBKYR6Ht9gvIfbhuKtizoyWbH9YhaV8ZIsbZgCC0bbKc34J67Hw1FeOMi2kilvLCIMtDKGzDIYMXjnAKmJ6ZvhXhehoq4+5mJaJLsQncjE/sPlE1GewoVDdFSVCljGP1dPlUQPYlRg0JrJGSrZTGxONsTI5+A0s4E0lQmKVlL5F2TX5Q0eApawnW0Jp64pl1hkEDcmWywnWyHxLsXngzAMOzeihZbIZGrsdZwFiBv1PAuw6KtkISlNYPaeGRDIiQm+h90xEtYZNEMly4O+LYsDQU4SENEDJKwjQwy3BfCViOpDSQQeopK2BCVDXkOolYuaSImBLoegpKF5oZeXRdoZ5lFxkHoKSjYWi98mwwYWiMg8sSRPBKCf0Ca6FrWM4o9mLxO2L0wsDhUnNTZrJEQc6NDrFF0WGxqg/qIieBmlMl7LwwrV145ZpVZEyHOW0lRLS8Ud6FoOMFFDw7ojpw600hsEIhqqDGkVRtcK2IXmnsYR0bRTlnvii63HkjsURRa9w16hK1jBGKY/3CSYotFF+dkA9G1ZG7h4Y3uwdFWT7cJYg2rgS3pZDKo9hXUUohiCFljG9FEOCvh1eBPjfCjjwzM4M9kjFWMSzNjwIe0UvjjJNDWtClghl+gPKjLj9UicVnZmzrWIRy9YnMIb2SDcyy2ghlox4azI/gNBN8aWR5xaVy31w0dgPbsbbEpw/AZi3fgkrwh4l+RORWXxyr7hzX9CsISZsd2wIOCC1rHWuvgwyoZBi3G+Oywdwaf2JJKISKs5wLyzV+QQq0cJYxjGFzLxbltiRUvXCVP1ha+R5RCFylTO0WeVJX4I/vGRv1zGbF/ghDXKsgnWhSk41m1owWy5aqjHP1mMmLIHtT7PmiG4McExJUPUehvIQlauKLID24wE/Ao6H4F4PDFz0+RtTaEsZt0xMCaeuUMQS1IxPwJm7J63UJ8D4pslke7o/BqMUD2BNPReESQPc0H2rA2xnySUvCOwKxp7wLRRWxcNiOeMBtTrE79GdPRTBDLEiwQsBtzh3CNTLhmWqW6Erw0RWx9lwS7mxxr5ELEjeeNZG+BRl2OI3WJrUiE+zoaN8JSsjcZ5H7Yp3rjV8ifD26e2JSDWSiY+MBMsRU98KM1G9nxaYYLAmKn5Cp8JfhN54alL7pjwyt8Q680kmsjLNDezPGX2cVGQtCjNhDQvkw/sNZ/wAFmynop7CHAJYtEia0XyK+x7EwDRbE9CPYDH6hsugySoQA1/0Mo00j7Ab001Tp0IPHBKpo2bQxGLw+F4FPbEsaKzzQ7BMJdi3MoUtTG0JN6RL8hFGhBnRzEFrUTZgJp5GiEz0LcetFVXqE74RimU6uE2W6yJ3sS0DI7W9FAIVWcmhZgSb0hL2KaRgZhCI0obvQmzDwxxpiTjZJZcE3ENhxPE4Jsw9jUVJwUbZg3AHNxPFHQiIOrNGh4MJWHdQsJBEK2JlPRLcimtRDaK9DvFH5PCFEDYhq9D0bsYd4yRpC95gWuNFZfI13gP8AtEzMvIpA2CIoNmzDYomuVsCjpLT4aT2W5GO3XfKKhOU7MUPsRPZUNPBkyiGiMWGr8Si0NmE2xY0ISsPIxMslKQu1/hKNuKSQ+3F3QMdKFIZ5CNo3whYxmLTK+gZPAih9LHQouTSSP4Sw5dSNDF2ei4xxTZ1iyIYlnYlqWSnsZc0TajJR/Ri8kVTCFFLylwKJvOGTAZV4FceGW5KIoliHcTjAtFlCnOC0pWMa14X+CCgeBotZG2OIhhHnWiKiDojYo4wCyxcrxHS1jOmBAHwS4RhkxMU/Aq7RXnoSZyxjYkYJOVZftfOLIQ1JEWiEPbYxL7WG0ssedY1zrjRRcP8AIClztiyeQBHAV7R8QcktrIOLLEtYbecJs8Gsc4CdjSSOuMh5+A8+K8NWI3nCNCVjFp7GI3guS4R0PMoLLdDIkbaY+b9coUathg3tFFAOfsWua+BDEh79AlSoRtM/SJlvO9iL2CVaFudiKBns8hCX4IJC6CxWQndoTVvg41GdSsbxMIWKuRNGUaVi5prWR7tRMyGy9RoYMTTVXFExpYMa0NRJ6GTYhI4k/Wv8HNhdxCTWmWjIKksFMl2JGhS1iUVBCwpWbDnWRnLEIKcs7iBCxp4I9gxksKDoSpBo1s8aXkWa3B4ekAtqtOriGhrdovPbIRu+h79B6iNwSqF0cpWLbPf2M3noQbSU9Z5AKwCd1wtzdDnfjPuIZgSGrCwZaZhPJjhD3wl+iMsvgb5Y7CdbvoWssXMeGIWU5q3oQbfkLYcL0ZGmBOjRGNR+GiK2IXRkbGL/AAmUW6MZPyJ1XisDG8mYwNK5LAdfJGtyE+xcNNhL0ooCH+oSEYQtWApZufpGy+OH1yYm2fgpy441u7RML9MVbr4LrhSsChOvLEd7GTSEMJUUDR+BLaWLOuGi2LwCFEiM3piuJizVF6uidB8bRZYqz+hFItGcWx2kx3DAhwzA+E2CRPYxqjV6PvEhNxDO6Rn2WYWkMZ4GmQww+EpkQu1jpPM3IlhSgxbs8glmPY0SstgxcyCdypLJSSxDGMGN8llCQXCtqQlf7i3PL45RIuDTca9qMVoxBYTBI9JMLCLBrlpl/wDILoduHyKkloq6ka0UjeDK0wQhmOxJtJaDjREsBIq544buC0UK9GMs23nhCYjKP/0GWXDnZHpoREbrwTtiOgkVQ8dw8laF3pFfVCS0Eyohsvgchizka8DTw9jZW0J3n9S9CLZdGhqEFXXY4yMAX3MxqJy2xviIZFA6QyIwS4jTK3EIkiRSjEDi7Q77gS6XwDS+ORdnpeuVkDOyiDxsv/sagF47mh2NlKNJIZQOqsMcQ6ZVG2RChBSlpvAqkPGS4hqsIVK/oXERSlKKZvCMaD8BtmRIThBGN1WmQrJFdxJLFwbb4SE4STrK7AYRYRkJEI4kMMLIkVZMQ8/yKoGs6GkQQvYUb4QlaFgkQvqKslX0amaUKLIixB4ThiEgxzZlusUlMClgZeK67Zk0yxC0blEYjbrM29sbHwz7hjwnjhDX5EYdHIrHwmK6+PhqiNspM/8AZ1wmQFei3hCRBrNHJ/8AZgvAxjQjSjw9l+HUGnhwTqqLCZ20FvFKK9w1pwwVSFYjLo6Zb8ELGO8EdWtjWT87I9dDE7nlMpksGOohuhu6Iy+OMTvFKUWROFvyCFScfocU7nmiY4x7hGJsPyPIxTwxOl4oz8K/wtMsSEhxwtm0Pbrwa0fBsSJOMN6A8A5PIZ/JlSHRkSIKaxzFgQxbMgGnolA2NiEhRWQugp48ZifRCDcSGxCELQeQ9BaAqnZkA55CIQ2UQ2kqxHdpaEdIsjSLY/8AQkQLjA+EZL1hDcJSbO8/7NSv9m8D53b4vDiI2/8Ao+n/AOWIa52Iapy0TLJQnYpP/sxT0yHoZNCmDYbXwdI0y+WWjoNW4xAO96LzROvK7GPGuICpUYV4fANO5QzInByZ0KYnA1iQ8YCItyP96E5NzRMdC2RhpNf4YdMiMgEpV8KU84FImK4oNKb8EHBC1c0o8inEsMYsnke0KULtdD3Fv7a/wQbS1mYkWeh0MimrGl7D2MjYgkNpKxDQPj/tKov9iuyxo+hm8wZbxDQus6FNsV0yaRkWz0rFeHhlEqJQW1jN74EEaJCYe0SFNayQen10LV3whtJU6zBVAUf3Dg3/AAVRL+hVJkbl+ongh7LaxaEGtw+eGOvWSy/8RKn2Nnv6iNOK7HKT2xplke3oaOhCu/8ARTVCc3saeuUJrJcLh8a2RvZgP/zBb/8Ap/yoix9mQndcNWuHlFsXZi7fnZjP/wAiL/jGXgij0MmqhpX6FG4PB/YQkQiyGif/AGZLZJ2qZdmUUm5CqIo4VZH6L/SMEKXsIOFFKMd4UpvK8jGoW8IyY3PXwLWBLrI54f0fYHcCHZoWlQs8JwWxl7Ci6IMvK+w0n/wj+7Cap8fcWR57GXbGNmgFxuaRNMh9BJkt1wqVtApffDSexFUQuA9A6p8L/CDA5DEaU/AEloN8GluNgShoU8KOsozoIYheCLFjT9XkSG0tlkfFkJf9wzzoSxDfBpuNvH9hCUi2S6RznQhaHs/0ISvY3w+6lbz9uGv09kPQWlcSS1BQgDZRGuxrAp7Cb2sS2YQ1RQbIYt0glEMS3Vsy6Hwha8h3Zs28j0f/AIESV/8ABm7X+GnDp0LOtmweUEELpr/KJ5rX9Ctr/wCDOkylsU2PD4FeOgklooxmCbiNPv8AoZ98Tsbkc1LDQtDCTz0NaKPKNaNP/jMoyjY3MpOge/RdVZEzf0lKU9qGv+Ua/wCUuBh2I9SIwyZJ7GNiExBAwzoaTwx7dPArsvwJY2S2hSGylGk1kRkHmwRtcVG0xVibwwXkRYil4pl2hqTTShZPg6uIV1whRIil4Tg0kj4qB+FwBJ3YlFgo2NlFRPyOHHgeq6G5g9IhnpksGLwhNNQWP/8ACCbY3s4mtL/Cn/pEiRDY2b4RJGJoCsit6GVRNaX+DFJf4KfY2XlhqaGRiG4dFE7M3li+8bZ6QosDGxCJgy6cMQsvPHQF937Mnf7GJn7HjiiMGVj+wvQeEWWJbs/srp/Y5rX9iGIVIUVR5ElJcIwsGIp/bMOl+2XQhjYEpXtCU1SHoombnDU2kPnSHLqRKfGwRtlh6G78E6MltH/g3/yEEFNBLUrr2PPKZvZ/8MP/AIg0dDn62MvIeK32Wqril4WsY+uX4EP+jsQLUlGTn+SHlc3lLNGE6EnRnrwQSS0KtFL8MCXJOEq0LIeOMQEXim+FVvEX+CKJCjZS3XCQ9ge8IfaUhgyCCSTBS8ylS2PjWjBFk2ERSGVezQ2N8JU0uBldZCLT+xQxrRL+xdhZGy8qDXnz2MDyt0M9gIvRgEkQQUb4Q5LvZ7IawS9ig0El6EwkyJJIhujEXp2Tw3BKPIib/wDhCdqfoUkl/wCOHw9MkBkuEPJ/6G6//g25M/oZqc/oZqxsDSPlHR5jArvWIm6NTPRmWCWm0Q+F57lRt7KH9Yzb0LbocvevghqqMa+Vr7lPj6AJWdBp0Cd4bc4o1EYxYMDZPK/s13/pCY/kY0FNy+FKISBGkTeCf2LbqiX3O9CRiKXilESRkVUlEKEVyG4MToUpSn9Nf4NjZeIilXkVgGbdHcSonsWUQ4cGxsvEirEzFMeRaymi3EElLAuwGxsvCQl4MDY92DLdox6GvIJhqC4G+NiwSdxDLy2JLVoZQ/6J/wAgt7/oSE9H2XA3wiwwrIQlZu40bBYJNYz+hHct/oc5sJXA+FT1BDZKqbHLYEKZO4PPQuLISsqVidYDZaOtjRI6yIy0G9rXg0Yf7GzeE/2NkL+ybqHzgeWI3XgTEIZ7C+Hm+xbRa9kHr+yk/wDkPXcYz/UsihkdOURxsZT2KaqSn3Gnr9mHgYtsinHp64DKm+K5KLriEXox6LqyEtoMyhOlM8scvPJpArqn6IZk14HuSwvHAC8Xii/vFhNbGtsfY6mn4MIciWPJQSdWBMpSjRKyjo6X/sT4BCTL8DbJFClKx/XgRYKh/wBa/wAGb0a2JKh7dWf8CdbVsit5NnIahESg3f8AYNlNiXkaNY6mYGiFW0rN/wBEhUWDY0Liot4S4Wnezy4/Cv8AQn9/0SCb/QuQvNYaGt9gxEhpEK8q6/I1Hs7YnyI/Yk/YxvIYkY2/+GC1YFwxaLAkhLwNE9C6LqcCT8P9ibw/2XiOv2L15Y5vs/3lPCpuVsbirEz9BTJ0KcL+x/zMSEf2MK2mPY0moJzHBq6CYI0M4DEAozj9kKOL9jSe0v2I6X7DJqUGmVkhqiEIyRsSIMLKX5FIYz4ELYaXoQ8ppC0rZDGN8W5CVJxoLZDL2NJGmVnk6ESe1+jHlfocfa/QlkwyS/sHxbwNVVzl4gpgtC1gdBv+i+/6L7/odLZJMY/0IWesTNaKNmBJLAhEtMkG/wChrVP+hMzZ+xlYpQ8bPtxpLbPYuVZvGN0D/RgBv8HgwZtvjGyiErHN19IbvNlTENg0PXlIIT5Jf2UZ4CSrJhCylsTf0RzmzRRMwkY02j0R0SQrFD84VhDnhmMImxK+WUvDa0ErlC9lSVJAyRY87hH7HNMipIomLT2Ve0SJqlTNydIt7Cjpi9GfY/2Ng059xEsFN7Gm+Ao8o1mxWobHDdhyhen9lf8AYtv+x0GELBSrjZodjFK2xJK0E9Qo1m0j0L9kFr9hauIVXhfgZKxmW/sGsI1DZv3CEiMHBRMKoNuiPIbJVfgeBj/1CM0TZCbBK17Ex5wOlHGPQp1UvwZNP0N+n6M6exKwtdpRcI2EmXsojQ7HStn4H/wQ3/wjB1f0LsI/E8ll6+K/5ZKkouVMQ+xv0X2/Rfb9GDs6Z552FrNWJ0bbfvYiWC8poHkbYma1jIjumTClyW5Pyz3Bl+C0jMkzYp4VsmtpGo9nUySvQx+vpcKXhCJIxrgrIWqM9BJyeYv8OsKSsZBG2DNtgRgilKUThEtGXbaGPCL4CG4ZhWMybaFLFxSlGyf5EIarwRQnYIZvGYT0xkI0KkhsZRBKRjiNfXsyJkzEssOvKZF6MTf9hjYb9mBDHwvDFQ9Pgd6Ah36soNDTatL9i9X7E/h+zoJJmVLLGxlIKtiaK1CbURD0W2SuxFHpD2wLaaGC0vwMyo0lCG+eh/YIQkQhMpieWRVNjzbX5MQaFX44WH9Ixq1WWJXOx5Qnw9NNH4GNNVYFXUfoFZOBSUJatodUfE2I07GPyJi4fM8Moj/qNP8AqNAqw3+mN0rEUW9f2XpFEXjDJw2Dfofu/RPl+hql+RK152GzpxAFLymISMZiaErsWzOj8AxLItZ54W8Xin3E4meeg2lQqCIrBlKUT4omKc8b39hCuhLiQkYELXO+Wy8rOCXA4UsuGxJslGCUL8UQDrKbDJo/IgsiUiGy8qmSYKZaQn1BThLwYm8MTvpkvcPHwQxJvZiJnyMoaGzaQnCI3vD7kJFhCRQYzZYrHrf2P08HYzxdiZ9Ieel+xuVJCCppEJNDFiKYAbbfAmIfSEzZhMkG9Tx+R+6Ei6hjHLGxZ2hSUhpzi0ePyLZVO+CTyg1Og0vKFqsxoJW9LHpPah5WBMohTExtGzjRguBjMWGL4IQGtHwKJkeHGZGn/UbGbsZIbcM85R0KF2LeLwmNXBOqEWqJK5F4TbYzyXAq7KUReZAZXJCOURgYEx+wh5ReKJiE2isRSbpC1mhjzkKJRDdKUb5nZLCG23SqzBii/qNkwiFvDZRs3wq0JXOy2dDbSHT1sWWGPbDC1i4vG+EpokWglLpQtsWCTwxJd0S9hb7cNj5Q4Mfu6PvB95EzpiS8hL7iUpNMylZY2XjJjG6RCBpMa4Y7nlBjM/8A7NH4osP/AHJMaGzBBulFiGq1FjDEOoGVuC5p+xjmLJNBiHBtDTBotqGaTQmLMiEhqV+xkpL7CipB+JD8CEl4GSQRXtGAmnsaaGUQmRaX8itmqD9kV5RH5QqpkmHTHTbITio0XiiyPXSPpAvQVkkHsNUI80HNENUJ8UvGDaYO0GsMxgmnlxT2JvjPNKPJXWDf/wAAu7iVXQJk8CXv4XjAxhpSI0rijZSiV2JXIaLQ8JJvIzyZDb6GcBC1iKN8XjeCMGLTA0brmtUbFaGfEU0qGauDZTZ9xJrQ/CuNjYm2hTcJTRTRdiOQbQx8qCLAmVsErWTa2fcyHYVwaDtwtX4hjZRCpT9FtEcW2JEth2G0xPAInQVNVG0NploPsf8A6HGqhPCNC2IV7ELWsaIfsTDad/kXlEzNjS3JDpGSBibbxkyMYa0IyQnFkts6wO/UVZ7a65YorSk2fgLTD3GxvijRKxiN9jKgQ6j8U9Ad4MCssRk9dejQ4J/BMd7GQJqmz1j0CI9I1kkLiFQnNhmsfC8fcho2bYwiIZ1wY7AhLeR0NKeoNoW1+NG0lWUx9BF10JOEIadYeRrsdgUzXDLvtR9uKSfUV/RU1UUbKUaSVjbUXYpsiQ22GhQqaTLGiMNtZEp7GvD2hspTAk+itbO6GL7B3DUjdBeAMKiCpYkExdPY34KZFkXseGFJ3sbbVk9Cegl6jzEJ1VkYn3IRRD4QvdGJtLm2eQhncFfofaPXMlVmSOiFjGPyIYg8KsuNdpFGXkXYV4FwFNMFDdgLpEsioRZdv6F6GZt5EWZEy9LRHTwdETinuQXf3PJD+Qa5hqrYiKmDjEkgIwTxS2InB2HGdRs6A9gfsxG8jYOx+QiGnYvYjs3JaRRLSKi7kngyeDGvFjCwfHLa7Lx2K8QuVrTL2MeTHmJ5hryCW1EEb0yxQRTs1h80aJQ1v1jYmiiYZkBT0JvaODK7LTEL7M98U2dDTY3MIpl2sjZxhniO0MveY7pP7HtVCBUPhfhf4S3t/XFFXoSIMstfLsggS1kaSYTnWISIomMfkQoVF4WcCFiIoK8jDyZX8n5mfyJEiOzajFWvXQyNZQkmONYrxkJuHgS6MewLyRM7iK0MghW86eyp5XCS2MuiQid6EYoqFwqcTzxUWrELcFPIhlmhDlirEkuBL7C/sZpkF4Ym9TwBFYEQ2SeM0ELAz9WUvPDuD8iJIMqw/IirQXoETrf64ljLGDraGqUR9R3/AOx600K1QhmNrFJB6FR5L8iK0gO8oS9i+MfoH6CRRGNbiKJwyrcxUg8h5UZG2YivKjfhG/CNs7wybTQ2mPQtaPuVJViV+gtEYaGnWNoNoKHULIFQ2ERDZnhZMh0/tjFEISMdm3g0acV2xgHRX1MiovhlNjm7+/XAB8UcajNoDfLGODXJ0OjsXE36V/g0kjKevwNTLOhC1rGhNV7NBBt+YboSiiHymWfuN5Qk1s6RbEw15NWD3QS8Q662oa4pRUi3kQk0Vd8VbGxVKBU5KDyLQhsThbgro09eiCUohsSb5CUK/uIuuCn5xuzFqrO1hTJ0oj/dEAODwHGISIpTi+Q9gdO/9jK7Y17pBMv7Fbib/sWEU1G0QZ2iKaIIst6IoJGuW/sLDb+xYb/2PzJ4J5v7F8g+9j1IImoxszXQq0C1ol5HwhlWgrrcnup5ka8w15jCdQnMTN0xlBMMW5hnsZaZqoTMVAsmKPMiEQnC4pINCfdDk9AWS41p/Y2Jl4QkDXRaH6SGm6mUUtES9CqJi3B39wRLBaXhMaTUYg6gi9B9oYeUIh7EqS2NVZs2m2Nl5TKJTGx6cC45hrdHc4P+tf4JiWM2ILJfEKdEZ1R5EmZ7svN4oyMj8MY8IUsWzElQ68h9wXuM84EJFxeKNRrm9GcWBNQbduxJJQYK46kghIkHxRoIRsMfv69j9A3oSjXKMjbqk8ZPCQY7I9SoemIxs0KbwNh2/oWVnoi7Ga2M60kfaheqRj0h5JVE5yg1azhlgjf943UI/LYhGVWkekJ4x9IpPGJGh4Md7usZp9isNRjt8OuEIV+wmsjNZztqeDIvQaCbyBatCSn49jpvS/sbFw1UE6K6J4Y05XAw0InsqnaxVWyLUTbsREPIuKIrIU0aQ2vOJ6HFVq6Oehjd7iMOaMXhc7GKjaGl7CTphq2oY9RbLHrQhCl4pSlEECeKPddicZRsPwv8PANjcNz4fRRrnQtIuaN8rI0XI4PQzbFBD2ngYwrYFjReaSmhz9zDNmO3IzTqEwUUxVkRZJqXhsWXxhkYusIdt7QyxhCC8KhaGlo7OGh5cHxYhTSRj7AEqhbGyl9wR9sJRsKypsi6c0Do2MbhcSFS3oxrEIpA2spi70/7HEJODnj9A/M/Q0nYsJINpbGxjIg1G60JYnw1VBNlbITpIoyzGrv+ieUgIUgxUVGqRKM3paZXaEnkWSTAhTGETTXofgIEfRYmnRS9CHkL7At0eyl5QRoeQPhiruhISVE6UJ98F+ecTJigosoRtxGhFE/AjBjc4vwTKIqtjXAsZL0hsbekURhl0JXhMWoCwovgzQxZEaj8mZeRvsxKcF7CPehJJFzeIzAbbGWmx2xo10hJJ6E+BWe51k+GU3oqDD0i7Mh2yO0yM2tDopAkCitgzjhjZ5jFbPuJtGENYHpEGh6pFEFB8AR0Dozqh+IMPQNjrGl2K4JkSCZguKZBGkZ4n7G8UJ+CGtyr0XwQ3gjywzFI0WR6LEYh0yJnoJtbIHqMoZi1BtMKOvgbyQ/dGPLGtuJnzbRMYiCbQ7dQhwvzjSskNdlGiVELeaYyVEQasyVGT0xMi+C8IQ+DRjaMwZLbsWJDIEFWWUKZibWBb4RSlFCKJwfwAGTwyu8iryuJYYptFhSl4TKJB9rH/QhJhzyg88lUiObayUvySFYIdDQ/V8FrhZhjMjXyYkg3I3K7GKiGnVwVhKehekqsw2Mb8H3PsQq7FTMIeLwIBPA/OJaZ4QpwhjqIXwWbFWSEGQajGM2LvkIdswC5hK0q6JIkZmLYMfC3DcOyFwCExwJeQLyv2KNkF/3Ty/74BE3UYyMAiS7sQhcLq8Q3bb9m1cDtt+zoOJ1CeYl0ZKoSWvJb8hF5WOoaREMJ9G2Pwb4EimnkappukKG7sNVeIaxymZ1sVHBcCrymZRMlETJCZEx6vyU4cAaK+GFKNG7UcPCaKii4vFKUXTwRR5KD6wNssQkL8LykzqQ3RM5EZ2KHxhN0EmmGi8rJeKNIIbo2NBpN55is7LbBUpGUolXxR3o1cZEyJid1CB5AhdkLyRlVKQyPJpQfDGGu0UpBCw9imsxsVifdMT8GNGh2WmBpVf6f8SYzT0LVR8ZEkqJimgiV5BqP8QXS36F5f6GxTJaf9D839HkyPIEGqwtyjSELBRhcLYw1Sy6b/oQkahGCVCP+ojgIl6AaJkVgkVFWZDhCJENbGhBW8mM75T7WmanKNcqMqfkWCZs0J8OFCX+hwHwu8KQiFSxNfeVGEaH64vNIlEdoaTaRqkhHpDcnsysCbWRKUJGy8aGpxSlFbxCGcMZbIz31zS8SlW8sSHsxMtyDb6LkLWtjfAyg+8ies9FKNkvLCSijZbErSI8obdSPTwF38N0ilGbtuv8ABjLwaKbI6yWaJsd6gpq5foX/AF4nJ2PwVbIe2mU+3tDfDHGO4vQsXo9YWh5kyhcBkeAsxr8SHiYWTY7d0a+3NEaUuIWhCNuh3cMtNKmLxReKMYCRkwh6g/GGMNB53B2zbaGs0yGw/YXGKmlsU0EZIZJBMTCieCPJCd4RPAlywLt5b7KERrExcIxfzCDrMsotE+MmTaBCoGJV08MaQTohql41GuyNFuWBrzR7ke0ZuA/TRB1IdUmVBsKYuLxSiuTXY30h2ag2BS9DbBy2OoQlA0VfRiHIkLxRanQ0wpLVtCpVDfFEqNUiMu3hCO7R6REsqOA0YkKtBJWsicMQSZ2UlNLhRKH06Qw5lFaHXxAIWmyMGI+wQmpBJkY6bIDQw3b2ZRD0CAhN0QV0gpIyJMFBD0WxCoOGVPIVHewyV2y0ncLYoJegnRoS8kYdoaudHrHqEF5lewhSoNiNo0yqhGj0tnaCEv8ApC/6Yrl0Nrq4Rh7oTqBi8yEiJoSiEcG6+FNYbfZ7HlRHsiCGgT8nibDcNkZzqMknRAoBk9CKKYw1HvZSaHriSW5WPi3rWIajqYizoeHEJ8NTIl7DrNvY2U308GGixkMk7FJ2IQrcdYmtBovGe7Njt7GEz3wcxj3CdmN8BxkX7B/YrRiDoY+yNFJUfC/zjriTN0x4GxVlnSi8KvBKQIjCvgm7oviK9IenkaKJjzXXfCwMWFWXHwghSLuG0TyEvInmLzC7rYG88JEP87/SmzDDGVlGJk+wT6inAIiAxotXRMImbhF46GmUbIieDOF0WbbbH2UcdNLegndzvjHlJJdz2RIo+GvWYyiO6GWBnB+bb2bEyj/2P+Jid/8AQlrVfkZHH8n/ACMf/aFf/sV2hmZPVjVNCHoxD+y/1zlHj+5f/wCyGKuyb9n/AGQ+BmvTHLY12IzaGOhm0E+Psy2N8NRGU/ETXJghzUtjltaFpUZEbwLSv/oMJNCYhOgzbfGfkJdio8sXRxfrI7R2oT2IbDei0NymIohu+GX3/QxRL+hwjRUWxKIajGhGfo0J8djSixlbERLLKYHGeKa8kBsI7Y77PYYJMYuWeUWCJIyx7FobF5ZV8Q/E42K44pcaJhb0dMrwuKyi2Jj63IdRt1jyFuRNCFCi4CUpSkZaCEa0J6OIGyi2MNae5Dc2T56GUTwtmKDChCQOx/cX/ZEWV+RNsfc/5GK+Vf3FhcYE221sRq7XAtnS/wBETVE7iXoL7RJdxPeJ6DXATV1DdRogxtFdNBtmbN7svCKoi8IplcjgeDwf6H4h+E9Y/AJGCtPuhYZClqMz30Y3svNk0OuQ6nBPkAJOh5AnmaVDwP7hiVqU3gaoTEkTA6gppgdEMHUxBjoZkhkuNjcbH/ggIJdH34paYayKslRiUo00500G0EEE6KNcDfqQm0xPAiiJ5Bj2NwiiJoeqYIDeFwmRRus0N8UpRjXYuMVwiKGFYvFGRAkIDCIKcPPCUPBRMcroEZaCXIZPTvQ9bc9/KCEnPP8AYSFW17GkbAjGXhsoikfmL02BWe8VPJkD2J5C8ouxnbYvMhEXUWMn4F2t5pSdT2M1ps96YlSCHSZ6H/TH/Ihf9AUUy+xHJn7H/Aj/AIEN6/oNf/wKUDFL8MZjBPH0v9PXFJlZF/8AqPr/ANRB6D/65/0Z/wA6H/1xhbsC4m0L4tiWKofZkIXneyipGfdMalqZLQyUPfcTdOMSKvQrY+uhspRqodTyU0gZRo9J6uBuBDaDHopBMso9hKUoaLwmURFVo0vJS9FOK64MgWRSjfoRaxYQsjJ0NkygjbsY21zJjbEqUpsWBsonRClgSUyw6NsnuPaLzi8gvKY+NjLAkkg+cNRkZmBKBpdIayfGvKe88s7UFO5yyLXOC80cRoSusb4AS6GfB4EPbOzD7HCSK1/RPr+jCPLZLUHiRiSaMpidEOnNib/9BL/+Rf8AWG8L+hXLM/4Uf8qGS3CzQZggrWW0SL2Io8kEPA6pjFuTChDTDMassWzLct2YI5Bb0x2FvsgIJlIRDKhUG4QzShlfJfSNm6KA2muSsDFKJigmRtB7yyMI/wCnAnwGaDKNwTFAhBsTEuRJkfCc4OdbDKMICPt8K3RSmj7G4xGwxmnGj47GdhnXC2PfD4dD4HseuF8NHDbhjGI3Gr7Hfw6EdmiNAtIfwR/obOLbw98no0GguJb4ZobnabGhuFvl6XA+HvjaPZsjedTvkZsI1HQh64Yx8LVx6FoRsLQt/BmLfw6TY3OxbELY9iNuDaI0Gacbh7OjbmhbGPYuEbnY6iNWPj//xAAnEAEAAgEDAwQDAQEBAAAAAAABABEhMUFRYXGBEJGh8LHB0eHxIP/aAAgBAQABPxA2EIBFFsf9NP8ApIPT3kaf2I/6CNv78q/tiH9cf9/Lv7/7Gz9+fXv3LdPf/wBg/wDXKH7sobnfKePtdZ/q/wDY6v1u8v8ArfM0freZ9G/cA+l8y763zGjc+28S+18z6V+4/SvzPtX7iP2Pmfev3EftfM+8fufev3K/sfM+8fuP2j8z7x+4/QPzPoH7j9E/M+gfuCfQ+Y2fQ959Q/caPoe8D/D/AKT75+4/XPzLfufMp+58x++fmNd/c7yn7nzMP3PefXP3LfufMfvn5n3T9x+ufmfXP3H6Z+Zt5fpvPqn7n3z9x+yfmd3+28S+58zJo/TmWfe+ZV9T5n3z9xD7nzH6J+Z9E/cs+t8xt+h7z6h+5jv63ec/1Os+4fufUP3PqX7mP6XvPvX7hb9L3g59D3hf9L3n3D9z7h+5hx9LrC6vpd5n+l7y37HzCv6HvPuH7h9g/M+wfuU/S+YfdPzC/wCh7w+qfmfRP3Pon7n2T9xp+p7xL63zBg+p5iVav03n1z9w+ifmYTL9OY/VPzCv6nvAfufM+ufuc/3Os4fudY/XPzD75+Ycz9OYbn3OszfQ95V9D5n2D9z7B+5g+h7z6B+4fQPzPpH7hTf2O8y/Y94fWPzMv0PefUP3PuX7h9a/M+tfuD/Y+ZT9r5n1r9z71+4W/a94fQvzBPrfMfsn5gz9b3lf1vmWfe+YW/e94X49/Pr379Jij9/+y7++Yv2YvX3E/wCkh/tJ/wBLPreUYxXLOI5iYuoyo6ypUrHpU7ZliGM6yiao9pUTpK0lXKLiHWVKmUSNSr3iV6JepKqJDLKnVEuZxUrXaJpKjnESoiUygi9IGZVRJUyldJqlQMwCXGIXEz6aTVKraJZKiURqILKjGpWIkqaMC2JUognsStJUSyoBcSnpDmPadEBYFHWVFX0iTfSAdpRAz6KxiV3nL0BcoC2BiVvKm8q3SVxHX0NIGPQkCVCBEr0NYA4hQ9IBElQ9HMrSVRHOSO0DMxLyTMCVWYEC4OCDmBmBfoGJtFCmBfovu7otcxi0ZJrUdYxLiQHWP/gIHvBSK3mJ6LmaSoFEpiRxKxKufmVHWUES4mekTEcNZVYmnoWTMDpElEcErPSJiVNGMTI5YeglzVK1xE6TSVHM0JWZRxGrjnWVn0VOZVk0xmazzcTMQms1gRJTxGonSXKxK0m8q6qVgmbjg6xImdID2gWyqv8A8OsYAwY6yvMC2VUpJWJ+oTEOukKdJuYFsYpI2bTUgZlTSczWDKm8InpWT0GsDMqJUCuk01lawlM25mrN4m0D07SoGSFhKxDQhNWfUuvQoLtLi+7umvMYaWYIMzVjjO0ajr0jKlOsrpG+0MaxpiKjQ8xJl6CMMJlHlCEqPzK0Y64lY9KgSrgp9FQJoiUSukDGkSJ6OyVnSGp2lVEjqlURLenoCbQj2SvTaVfWJKGJHYiFejp1jmUzMYjA9HWVKzAlRIFdpqgWECNSoysTQ0m8bm3MrpEtgSjX0CVmVTEg9Kp9AlQKKlX2lVpKYFsGZUCEqyZgayoR6QqrgTWBAp6RJ0lSvQzmc+gm8DXeVU6QGAaQJlz6jTEIGJWIdYJiGkIawd/Q/V3RKjbGMUlVEvmPEZtcqEWawuzoZVSaErmb4leqo3cbGZVjxKSVMo+z0MOsS5YROZkQKm8TEq4CSoxhKwSmVcqJiUnoj6GkqBnMSIw7RlUxyzMeYz8xy6yszR6ViJN5rn0r0cJWY2egyrmhNEzcpJRAlbSqJ+JXpqlMq4wE4m8ZUqVAuFoawJpKWGP/AAvMMep6kIYwmITv6ZmfUKJVTJBuGsKmk3hiOsu6IbQ1gMMMC0MEuHWFGIYg9A9PpeWKpHSVUxKTPpozWVEjmMyZVRilRJh1iNHmJKDEQlSzvCo5YhcqNYlRnTeJKjidZVxzKlOIhKFlVMysymGcxJUTM2gYj6O8HErWMrGZiXiYms3iZxAjgmUSpt19NTeViOtTSVh9Nb9ExHvC8+jEm8rmYlyswL2mk0r0DmYgX6VeYA94b+laQNqgVNYlwIHtAIBcO0THoX0SVKqEqVUPQBhrAhpLgJqxYXM1cGVfeVmJn1DMqmZgXAYQYqBkhFhkIYlQPQaqBcMei6lz7XlEgblZzEz6VEplY6yokcMSEBZPl6RvqOriJRKz1iaRCokD2lT5SrmWdZ2SumsqokQlESZSpiVcSOEqGGa6wI6dYX3iemJWcR4ZUcsTMXWMYej6NEdYs8zaLj1rEqVE1l1GbESGZUrFSk1jpAzAmxKmkH01niBiBAmGUyuZvKvpKB6EVUOYF5gQJWZqxOJvLgRNZtKuMCV3iF+lL0mnorHoqViJTC0D0C3pA4jl1lEdZWMT8zSVR6JA0zK4zC4EoqBmb+hp1h19AtmaxCV1Z9byjrHrHJ6ViM01jXn0d4rtAuCl9o4xM1ukHEaxFmsDOY5mTSbymJifmb+jEIIhKlMzGyPKVtKjcISVKxLxHEvmVU/ETzDBe8yYGYusrrE1nTpEm8qOuJ2i2Rnj0/MqyV6VKr0dIkN5rOfSjeVvMmK8xxBcCU1j0c4gUyphPz6bdfSsyukr0czeB6JzDZ6CFzrK3zUOZUSiEblTSOe0qiGkzAy3AogthNfTvHFTK6y6IazECad5rKlU5gQN95Uo9AGBD0ME17y6ms2IMIQgvpX2ofq7s1iTeBGJmJK3jT0YGYYQG4CcxUVAWtY5jAdY5RKjK8srMrMrPorMSJrmOZUS41Lt1malY9KlXrGbPTeJ6bSpppGc+jKz6UMTmJ1jRElR1idZoy8Ta42+msSs+rrKjKoxEuJiO0uXp6JUGURzHBCasIeIa+lO7ExKqB6EAgZlZlVpNdYegNw1lTpMiV6JH0yG4FYlSvECzMSprAhNZpFv0rN8+iswL1YFTEqEq4wJtPiUMqDEq/Q0N4FMzfSBbDHofEDMvMIcyzrF9/dl5j5mKi1L9E6zQmWVHWVUKgNyqhXSDTCZ1mN4xjAmkz2lHmJjEqvTWJmVGBrNY4fSpU29KgzO03jrVzRqL6LmPMcsur4nmXn0YqVGMdpWYgxK0gTNSsTNQD05nEckcelW6ysROZoRLlVUqOtMCGSEDM7JWIypRDHp19CbwiQzvC71meYXDWV7QIGYFwOZXER8Q10mt+lDOcSrYHpWJVzDSVj00lcwKl5mhK5gZ1jrcxU3lRKhgnSU05lsqFTXeBZBbzNJpVS8S7ITWaQ0hkqHHoOEmfpMfq5fRcTzmL6JccSoY3jOqOsDXMGLiYM80q4kuo5lTepV+lb+leipUrWJKajFX6Kr0dprHa46R4lXKxK5jwmE3jjEqolytZpGfn0qVEsjpMVrEphr6K2iYgPoSpUTNQiiYQLiRzEqVmVAxFhmVAz6FzSNkBqEqxlR6S8TPeaQLZlgSh9CBcC95tTAqMO/pt67elAxxCZgXiV6E+4l6elVKzrNYSpU2zpLLl46+neM0xPMIBdnpeOI6zeVmV6bQhXpdTrBs9K6z7Xlj3nEdfSpUQjN9fSonopAQRm5kh1h6LJQmsCtNZ1iXDSVuzXMq7lYYSplEmzNCVHvHUmRAjDMSoTVj3mhLiJHC5XWOJoxpYzmXKjSMrPoKzKIlZlMrE0r0q2bxNI6SoErM1ubSrnWaR9pS6MCod5vGV1hiGblVEtzGyKhFZlZl3cCaa+mkF1KId5Qkr3hp6BNvSjWXjn0FRlSopfpVemnoRJV6yoSsyvib4zLsZUqzMJtjMreBN5XE0QKmkzKwTrL5lwwQ0mzBqNZswwQVmeCfS8vS46ejBuCBKzE6+iHmU6BCZEzFjZpDdGZW0xo8etRuBmUO8dZVyrlTMSViax19EInpVxKlV6J1l1USVL5ikQlRLjjEqmUO8SpXvG2VcrMrEphEuOs1ldYxziVpE0gYmjCOsek1lUMqG8rM09SSq0hg6xNJrKzKt4leltR5lXNPTrLZrLmpBhmJcAhDDrPxNYEDGfWsT5ntLxKuYXDOs0WBcbuB6VUMymUF+gVZKiYmiAVN5vUqFIkqoGYY9d5dTTr6VDWaQ0gyr9WmPS3pD93diRjce/rVxlYlZ9GyYd5jbWZKrEbRaS9LKXK9DWOCBeYmZmURlR1iXEoqbStd/TViSsS7lZl36a7YjliJWJRBcqiViakqiV6K6RMys3tE9EqJMpK49KmUrPESVe8rrHM1ZUSVm/Q3lYiQXEqZhN5gQYgUwKlSsxJeZUqVmJUyZW003lZ9AtvSGN4QhAuVRNJtDJUyaTWY0mk5lWdYaRlVv6a6wzcME0bm8C98QJpNYnWUy7x6ayoMkrMN/TWF6VOkcSsyoemqVe0qbTX0M+gw0doYg5l44nh7TP6uUrrKqXbNGXe0MSrmhNcxqmGCpVkFw0HMB1uM6sFLN9JWXAlQKrmBZEjFXU0RjHWVqyprHB6PpivR6olRwndKpjakSeIm0KStHppHeVUQlRIFxJWJoxPROsXMGOsvENOfSqfTrElSsayrP8AwrFyvTL0IYSqITVhk+jlge8NZc56ypg0mhiMqmas2gYgQbiXKqaZly7qX6ViZraZ3lTaECpWceggX0gSrmSaQ1lZlHMPYlVPiZ0mnpXWHRl9fRhpLqvQ1g5nEuLNIYZrBqbQPQ5gW3Kg+vuyo67yrYm0pNpUrMqo6+mSZJQwz1lDpctAxHWAF06ypVTWJAr0Imv/AIJeZVxKZfo9pXaXc309N5VkSplOqJKuGsT0PaMGj1S5VMSN+iolxirjKohr1jrc26+gMdPWo9ZcrPJERiTeZQXAPSpXqFt3KlKwKlwbJVyrek2r0SBUSHooVc6kqyVTKx1heus3m01le8CVNZVxJU4lSoFkT03hO8C2VK8ypqhnaBAl8wm8qpTcdZZ6OdoHppBGHxMy4YIZmXp5J9vyzaayqzLxKlZjpAI6+lWeh8TeaD7y3JqaJnTkqVxKuVUqeJQyi440lYiSsSllMqVKqZXj0WrMqoteiswLj2nxKzEhhGKo9HLEzBmvQz6OGNbayq7xMRKjpElWzM1n5iVKlejmUk3lYuMq549DczEgehAzcS5VQIkqVrxA1lRMyqlQK3nQiSpvCVcAJvA9N/Ss16KlYlQlVcqMD1zNJWLhoeiZhibztAlVKzM3KgSssYrE3qpTWOdI5lQPSpW8SGJpNCDiXcDEJUqD6e7Ca8R2gVWI6MDHq6ypUdY4hmYA2l1pHaNZcylRlS71mrKfRImJtEqeIm/o8S629GVKj8+hKi9JWIBcTPEqpWLlUQKjmJcrMTMe3oIaTXaMqtY59FZiZlQLjKxAuVElROh6ksg4lQSsR09HLAxAxmUYiSumJripVQh6KC4vTEG9oErM1vaXEr1IboGZUNJUErrDMzdy4Yl2MqJiZhjaGYlyoZlTpAlaQ0jqSqjDWbsC2JTdTV4mkJeYsWtIS5bKgQJaBxK6QIdoG0SY4mrvDtAxNH0wb72zeBmBHMrpGZ9DWLKsZrKpjzEmE2GW46xUdSokqMoleiQqo6yyI6bejEzPErWVTEiTb0SoRyaSomJtE39HMdJV6elStZojWYk0jliRai+iVKxcrNysxgOnquVEIzmNXBbdZi5lZi3frVwlX2lTeVeJWpxAuJCcypU09HMNKm20rESpU/MqAzeVi4O1SswNol+hmBKm3oGYaemYEJhAuZJWYXGd4WyppGbgUr6uvowYt+iQxN4axMw9H03lVLLgSpcth+3uxoTAlUeiSqiWyojxKslRKlQ0xSKMWkNTAtQi0rECaGkc7RMxPRuBiJcTMSVU2qpmprH2lXK/8KfTaVZHEYQejiOsQjKY36Jcr0SDiVN/S8Tf0rEq9ZVHaVZKzHWLcd44TTaJcUbwIGJWZcCOWVTcO0r03jrAlNs01naHb0dYjWkqpUqiXWkr5gSqz6bypVSpxt6VK9fuIEYEuVKhhlXKlXK6SpXp4mvpWZVPqeiVEuDAzGEreVUZtAm2kS4cSpc+r5Z0lYgVKjx6JLqaytSVtKlRMTLmGpvGZogC4lelkdPV1qVKzKqVvEbiQqJHKJGURJXo4lTbrKiZiRMQMR0gRzKxpHMT0S/WpVEyZoysSmVXj0q5WfWqiYiRLjr6HFRqMTEBuG1ypVypUrpKliVUrHo6SuZUCrgVtK6RIayoXCVmBKlWxagXqTaoOPSrZtNllem0IEq2GIZiXKwQM+iYiaysSoEIqVmV0iQKmvqF+gXKqBUCFEdZlt6Eq4GIQ19O5h+3uytPTX0qJmOUqViaMdZUqBzFnMdE2gh1iakoamm0WpvXqmfQkqyVHiJG46zsjcqVTMoR49AzNXSawJm5USVKRhxiVj0omDiOukEqUCVe0qVpHWVmZSpgTaVAxK9WKr0T0EdYwSsaQz6Khhm/o3KojrE9AuVmBUqLNZVTX02msIFxKlY6zvKgyp4hKuLDfEMmkGjSJtAzKSq6wIErMIES2ASpXiViH/nWGJvNIGzCVDWPSEqaukrEriEqBKr1fS92VEIEDEC4xMWQMTVH0JA9AJUOITlhMFdzPEXEMPpvLiYlw0lXKxcSapgiXKuYIbyolPo+m04iUHpWYsSpVXNGI6vojHpE9K9oohrmLcT0rXmVmXUq/QlSukCpWIkrpEusRJVRJUStowymAwJWeJcC5Rc9iays1KWB0gawNYkI4MSpXoxxNar0CBcdYGYk0laRPS0BCIXNE0hrDO0wx6GJXHoSyVOkCVAz66+uIzBKgQIQ19K0gTWPaVmBAqaTUv0Lj6Nl91mDEqVKlRIkqA+iSqZ3jXoSqAcwqVLYSlJUr2lSsZlAR10xKAmpEam1SsR19E3hGNppO+Ykr/w5gSsyrglXyyomYlSm+kcejE4mfRVGkSWqIyrJVbSrlT3RNIZ2iSolSrzExKq5VxJXmVEBiQHNypV1cYqvRMcymfKVmVKlS61uLGbRWYlW4jL0mu3pUYKZVyq6yqZc1gYnMKr0C4aQN5q9CdICTeVcxKtlR9oTWUT8Tb0cRPSuvoBcSpo6QSoESY8w5hrBJUCvQISmD7e7EgS5tKjrKuUO0DeBzElTfiOes7wekcY5AXby9cS2VXpkYysyrZjSaE3jfac3NTEcwlcymJExKsmo2idIEolVGVCKz0iHE1xGVcSVZGpVypUekS5XoyoQUIFEq2NJUrESIyquOkSVccuk6SiuI6+ivaJ0lVtExKqoGbmifKJTDPeU3B6HXMC7ms1xpKhrN5U06+gSsdYEA0qBmJ0idIGJVMu5UrGYFQSwKhMyocegXKqVAqZWbczaVHEqu0SXiYS5VsqnE3lX6AOJqlYlTpKlSsSnaVzKlZzLPW+0+q5YwP8AxVyqIaejiNSpTHXHp4gZOYFIMtEYUYkqVbNErSJ6WR5mYlxisSoFxKjH0YlkMejKrOsdIF5iSsSqiZiRGcxJXoqVmJcS9vRg9axKtlYzK4lES46emiJxK9Ct8xzKzPxBghFff12m02lSm4a9Y6xJXSVR1mvrWZU1eJXocBK7+gWXvAqVcplX6DCbQGBAjAjCGsrM0lcTbX0qoeuqpXWOk2zFKnE3m3WBA9AMC8TiUxE0ibRolelUxpmjHr7z7bl9NJtMzRmVxKlZlzXaNetV/wCAIS8Q4Yjl0lDUqoStJT6VcqsSvTeXZKxEveMu8SvRIwBMVmVExMxJtHWOXSJWY6zX0E3iZiVKz6V66yiBKuYmKleh8TFysyokqVKlcEx9Qiuk1QyiBEgelEuV1hiXNIzQZWZpNCBx8+gRInECoFendKz6MIEAYHomJVTF+prGbenf1rErGZ0m8qOkqxlRIEqayrlQK9KJVzHEZVsqVHMpCXDtKplT7blniVcR7wyxcSpWZrAqOkOWPT0SOsrEZVRMgzALcTVVAQGYET3mtRG/SvTUgRMTaJczKzDGrEldJVwMSrxKSsxL9K9ElSsxfRLltpUq2Mr0S+kAnLaauk3gZhpAxKtiYlYjKlNxu4Wv0BOPRoXAxKxNGOYTf1rMaYFsdZphlRIw56ypZ1jlKmsIlwgLlV6BiVfoB7+gRMypVOCVzKuEVcqVZAx60RPQziGkrzKzEzExKwwK9KlT8wlXLzOIwa9KlVD4lZxGNSpvAfQX9bLGoETMCJUqBKDEzzH0aiV66SqmTEZexEqBaoj659dPSogMdaiQOJl6JcqrlZiXAlQmNJU3ieisxMSpz6VEslejSPeVWkT00SpRtOIlzR6KlUTRKLjExiVU3iEp9VZgg3AeYkpZUpxDKBK9oRCpTKiZlVGpjeJAzKziVKJWZUDT0DnSVE0iENZpn0D3lQgXHDK6+g0hiBcaGbSscwmkqV7wKlQIkrHolQPSpUC4xWIlQeYQLlT4m+sJWcaymJZNCas+lPM2H/szWZiX2lTVgVKrScSsxx6MfSq9dUNSJVjE74AUUKOOspppAiYlSpXSJvKxKrEcsqVG5q9FVKicRKD1VnWJmVEuPEqJRKxEmkZXWBmVn0DCNn0rf0qGWVNusTEq9okrESJccSj0MRG7EOZqm93NNJpKxGBKpjrNoUlTZ5neb4ZSyvSoGYBKuVmVmd0CVcqaeiq9KuBUrE0how9NfWtYQgYgSibf+DB1gR16+jn06QJXLEqGJa6+tZ6ejRJTMymF+gYlSpoTU9H13LKslQJQxM49NZWfR09EjPMq5U0xAJdqzKMqmEbXEaZYLWYlPq7Sh9PxElelXvKofVuMqiY5gXNJ5m/o+lx+IR1niJXohELiUS8QjmVoSiLiGus1YhU2q4NRcTFZhDKHeWvtCBG7bmZnrU2AiFKFVtoloRrADFRqDgOcEKApd48xGSGpkrxKB1l6Sw0fdwGo8AHUUqfF6JRSkSa9JtGrlXEzj0b+mJfpvKuBHEqVDSBiayqqeI9ZeKmkDEr0TGsDeGZUSJDDEm0MV6Bc00mpHBExAmnpfOJUN4E8w+YdYlRc+hKp9Al5g0zAlU+gI8TSIehW8SVD97diZmunpVTWVDE1iV6OfRX/AIqXUVOINmWBXaEsEShZnjSOhEohKlYZVxxGmI7+tR09NY5JUCMqViNXElRPSs+ia+iSsSpUTMrFSuPSus31mIAZQhPuMENKnMxbRDFgEDSFoLUQuqhoicHtQvdGRaDTNOh1is7wPdhtmMrdjp9+HA0/saxoq91/ybCV+eA5UGNTXZ3jEt+QPyeJdJlofkhoBSx2HWMGOkGEgbkBg9+IkI4AUjbJVrqpqR2w32hPuPG6W8UGF4E6Me8sm/obwL9EhpBNWsPQHqJvmVcD0JcqVAhgjuzEM36VAIM3xDSbxagYlRgXKgXAzOsrHoRblV6Ax6UPpWJV2QKmXWVpD0C2VtMw0h39D9TdlSmVExHBXrUZiJUD1S2VA5iXAqKo9FqiQ1pnKjs7TWVHLESiLUYmI+iZjmVK9KzEZX/isRJUauJUS/UlSnPoSVRHWKQAyhLtotQZbXI2X5RA2+qBMGbqqh5ibHbYCL4L3W/aXE9Umvu7RYawzVod+YDpB1Rr2TFguE3WEa0aDZ/TEVCtD4d4WNC2r+YoOkUv0tiYilKbbn2/MIRADARdqoK6H9WMcZXyTicVA/E/r3j5NNb1lAadE2dyY46vu/jDSmYP4ek0bEyiwcnSKt8n+Bz2lgL892SEQVmsMv5MV9ZvwzAILYp/2CrqOYPtAZFy0+Y4HUKx8kBkTn+0IETmx8RQpfH9pRmO4Mo7wC9ZghN5dwY4mLlXGpV+gKlf+GzWfSobyjmBZ6Gtzf0CVbKz6VNoONIHSVvCKO//AICV6srPpdPSOWBb63tLuYGJE6zEq/RfQ3Ya+i3EuOkTHrvMSsyvRv6V6Vz6a1GtoamYSTEMFGnMfJglYlX6IXHGIxAlRIm/o6Q9Kr01lTWOOsSyVGNLgVNZU+YLkHea83RmmZGj/pNM3kDG0P5t+WCMWm7GDy3NAfgiZgHh86sdKHH0e28GqjotPBA9PiM+CLijaXk7QyE4jl52lc9kNr1f6w8d3NJ35Y1AcRp1PEySXVmnQ4IqVDsnjvC+Ae68sVkWo/uo3i3eoS8st8Y5fL+JYNAFx2xu/vbmSLsTFebhF0CpfA/NPiWGOm+Q4Nl86QuQFI7wCjVr8uvEECcjULpAtew6HTh6RC54/kIDYxrWDkd43MPdMu3EtXPvnU/yVb7Hjs/2FTk9Rw/2Nu+wwPGjFNu4ce6giDznPswlKHfJ8OkrmeN79awN0Tlo8MaYniHxTHjfmzr5lC+vMmutHZ4NG/4MKsDlS5Tz6VmH/isQOsrtNpn0CVKrf0S4BUvtAg5lWZZgx02gVm4QzExrDEKiSolPSVNIlwNoErPqFSpUNYFQ59dDAuMt1g+huw9K6+malxcx/wDFV6MdYSpVxMSqjtMkYehCplDxKlZjE9KxEgUSqieYlxJUZ2lQlSoGY1MVAFoO8vuv0Qxy7uCyE6LDFiLyrPxBUPZAeWE7PdVV9jEVgG+hFXHzn+Rsy857bQVldXn2SnGps/ARwQ5cvZNUlplXtHS3efA/sVzcktmns9vLsf2MBGl5S+ZWQXalr2b943razlK6sqyq1tHQ5ZXZbyi1crG2g7Zf3wQ+DRqtV5esU6g/YX66wPKKi9WNNhdK9XwWy0EMPEuY27pcH5goKCGOCMA64vEvMbR8TUSOjmKlrYNyn5JYVTXU6kUP/BvIgdWt9x2TrGT4sOjm78keY2ojSPI7MtvJTYOh4fzMshqI0jyO01C6QGex+5ayaisnUYHYo/0DeU+sCMn8mrnG4P6ZrAuzkX5Jszla90wLL/Ed/E0kvNe8AcdwHgQDKe4fMFu+OT3NIrsM6e8sAYe2/cWBXCNfuZM07sfEoumsX5ljYM1ZPzGGk+h/cXBzlk9yOmQ7UPzBBH6D6KmhLzLzDFxLlQIFQyxgaSoHPoYIFsSiE1lZqEVCkCvWtfSsR1hMwygZiXKqBUr02hGoaYlSpWJTPoG7K9K9E6y5WY5nJK9HJNNPQHMrWBEr00lcQZxMHWFWVKjmItPXSOsD0rErrGJT6JcT0JUuDmAdYAtBwEZREYp/wJyp0aH8w17kj+Kh7QOxH9y0rru3sQpHq2PuwDi+9We+kD5DwZQZc2y29ggCh5TPsS5PpXwSiQ8SFjaD7G8H0D1H8v8AZ78fb71EtbXfX9jPZcbfY28xFV7iC/5FptVwHzv4lDWdBK7DaHg4SV/DrExFuJfe5/EFuWrQBEFbHGC/XyYeBqBVEVaZvp5D14IAr1tAruruzK/WKVpoHVYviYQyHYdCLRdkDFN6tU7+vY95Tp98wRKaEHAfyCU4gAAMsrxLs1bZnp3iiv8Af9jPQp8n7C/MGKxAlRwIu2/JZ7XFoBLEgDLd097JyRx9Nl4dk6tmA4BSo9BFIzx/Sxo2kTRjKjURx57PTSOFSURF4TaAlqzR7DeLe+oLt6O3ZlKgNSg8xLlLYQdzfxNNA5V2vyMdtO8vtq94M0BU+w6MQ7PwtXj+TdXWB5KuEW+ZRvqf2XfSdY/RUHjbdFeGcdcN/NQwpkbNfxcdjoQ0PDKJujQ+z/ZgnaI/pUXSHCrfcIrUpvq+IA0W37cUcZoVPuQMs0zN9koneAH4lQOCKvmAMrwsA6NwqHpfoaSpU0ZVwJmOAhriBesSpp6Vn0q5XX0N1BlQh7eh9TWVNsyoZQCMqV6fUcypWImPRL9QRcys+gcQiyr1lZ9ElejYgJANYzxMNVBXFQJWdJUrHolxLlSo6QNSB1gDjNguKEDEL+GAGCtdyz8VGFQ7U/khp32kSZi7rdl7pMMrwi/gIGLSaOPwERHeBg/E88RfkTDkHgK/EuE2br7FTTl1Q9quAZxwo/Fx1dzZfOIFYG2+gRRKrOVr+RbpnIR81nxHwoD/AEYTEHQzF6BBLftWn2NvMR2DWx/xEHDXp3dpgIGuc8+Zc0AdgJl3oJOezfvpAlnFqp1YMuJV5TgIg4DSzwPJ+IONPlCpLFvbynOvBLhqurK1VvWEIQFq7fMCPQHKvosvuHvMKxX3vBXFnZg38+IOVOsJldd22XW333i0manRBvwpd7Pv/sVsNx+6xgtqH2I5j0Kfesa2fBMb7Qw6fP8AsprhFOE94x6huss6a6rHapyr8f2VzUlnGtraccMABNaOhqi9YD8aARIyLsVbPe5+RHSEsQROYQqDFVvQbOkX+sEnlbPRmGiTQjF9DfFj8HZhJW0J4v3OwyYP9eZcwhtlO/8AEfUVs0+5UvHn4l/Z4mVdsETzWPMryWaAH3JcPSiPmqYLXbaZ+KZliuEK8JKPyi9kmjjrx/FxzwHFfyFx8C4H6phAvtipTY6l/Co57KHsJUADi/1QOuQfykXl0bf61F88csvyEA3St5fxmJgttV8MdpcH51SxCtW5FhHyH8SmH+FJUCnCB9mGWPzZCKlSqle/qKSqIZm2kCVxKidIFkcQZlXEqBHT0CX09KqVHKVKlZh2gEqV1n1HMC/TxOsSJZ6ExKlSvRJXrqiMqtIkrENSUErAxKDmaQNYqL0Zo+jpAGUIb7NEXQ60/jDWJbAMAzbdr4i9rmuXMqA6/CCUPUw792FL+B1hQ6qvfsRwshwCIm6zd+WGrJ6iv5AaP3j2IbwbKHvG+IPDL3YLcszkf3Cg0YJ/JOCuYfLGupxCrzcMC+3Q9tWZVvi/ZcDnBZD43lF74vFr94YTxZ40gwQLFquxB7ZxBXYvHmUMt0b90bFuZF4jra+C512eIMPwAz85gxwMAV6ucHVmnVbCeTl3xCwAqBwmJ+XQKPJsTKFmUK6BsRXD7EblgGgUbvPAggUc1HdK7s7A8QsmtpZ3C8urwd4VDIAAASgqmoZFIcIWXkDupfR+IrTr8Sq7RvOwj8sDv/SNYv5IZyM67IW8/JKaaRezAyvepbZT3JgYHuMOs9yUFFxgr+0+amPYyxZyPUlLA9kWcCU07Dh8mJX/AEAaRVAR1EZliRXeco7nPshF3sBGDjqkK/FHTcuv5NYZrrLAwNo3efRhV1GhlHSPkhEisskvONOHyVT5mgAdwle4eLJz3JYQGfddOvvCFYe68hqS/odyxEbJyF8beIrzcn5W5LquWE1F9sZ1fcakG4Xk/qPaEWDnCeSYXkp+TM0QXX+LJDm3dkfiOh3i/IlakcDLAPmYfaWGr2GH3P5GwM4P4o7fQkK8QHguHXuQcOyI/ESbeJf4Y26+VXvC6v8ALp8MPVxyfBlVfVxPtKI61/WkqBfml7krhB2L+cAITxMAFIyrJWIGYw0lWel+jrHNkCiVcqFmVxKzKlRLgYhAqVKzmVcrESyZ6+8H0N2GKhv6VK0iVElRIlMq5pEuUiXKgVG5UL49KzKLRm7SOjA5WXDX61P3FYuGs9/McuiUvyy3T7XP4g3f3YGvOZavOjh7EOIbqUCys6JKWG4S/dlS7Voy9orgepf7TL7uF92L8qyvxMFGdlXzR83AX3f5MpTkr8wJSpixfdYmooyqvd/krXIzfXzEwDrWnnSJtX1H3HHxNU8uL5jKR1FDu6EyfUd7rg+ZShyJ9xlZbYb8Gkp212Mh+D5jNe4sTyytELQHsAzALy9kWfg+Y8qPUVfLNhxFjnocy7gjeeLZ3faGq3ULumHgq1AE7rhtj7ZfmMA1TK/Kyj9rijBbDV4/4CZzBa1+V3ihv7kZoVbNdu9eD9Qm1ltqjVN2cle+PyZe6H9B7EfpyM7OU6rD7OXtagO2V5FIuyhZky17rKS21KXSEcIhN+Vtf5lnWFK0keoPct/cqQCaSBiog8pQ7D3Q6vYi3C1eWPp1fGw63L3p7cVyHtzOGEzT7Dluba8yoNFiBGak7FJVUkA6uLo0e83ll0seE2ekXy8IopKUPsanmGUaRQ/bc6mI3MvtI6rZaH7GpmY5sWj8C9mmW71EXr5lzj2H8xCpWhBO5r5Y6wSKLEBjniUL7mj5hgDOL3fzMLZhAWdzaL+Br5K18xUKd9qv0/EuBvHP9PEsvXz5IRTn/wCcGPiGwNXmdhiakp0pPuRtvXS+H+wRQP35n3JipegTyZmpodL99Zu49O9nMxEuhvvmHwKH5z8w0ScuPs/2J+WU+Ygo234BuF+Tvj/ZMa/NaPcuGX56ns3L3YDr3IqxuWr8Q3AOqBiVWlsfciN0m1E8NQ4hbFD71NOzdvQjuyg/qa5/DH4lfaOyB+YPYfIMK2m8YbUjwlMqEDMqpxfoZlR1lUSrl1iBH0r0x+xmbysx3lbzaV6s1SolRK/9EWoeYPdJxEuAJbJ+EYumAMUap0UXxFCi2AryxGmvUj2GJRby/wAxBEvA/uMHRxt9ogqkaOL5lJsvFqaim+g9pQlX4veUSk+bnsRDXoqj4ifZl0J8PSnxrNQ1b039idbO492IV9eLYLUE6j3YldD5z3YqKuY+IYZDf4XQhOpe49tINp2gz8E+sPsGscFf3Q/cwwDxUioh4Ws99E1KfgHZ1PxGJPS1xQwYsx0Ag/KNqqfj5Sxbtwu4sGr1tAJYuaGuOyv4m+VqTXZVeEtX3fEaM+yr7rWDqw+KaX3sZdWBMA/XSBP9RgBCLvtMUva/kekpcWgAPiW/5QUE7cH8+4N5YBznX6puy2z7Yl1SVnoHVihz5c5Pc3evaCMV7JbmEE3I4Qo+4+SBRIspAQV0BjGmEZ2CNv8AUtWfnKUtYrZafuLWJC/yxDbVF7ZNz0IEn1fMX9f7gn06FkiwzzB77dHw18nRI2/R+YIKbWBNxJaHq3Nm5en+IXo88jTu0Z29C37cX3lukYtvAvDKbOgd0D1MVz99zo4lv4Ydxj+B8S0ESSHDXWiOIPrh3W0dH3jjZbyuEyTAiKdt0VSTKLfd1KYVVcBufw7MoElkd84NlRfJFa1vCD+n4jiRdQ90OY14cVynNynxup8xMA6Dd5DHmChxqWGGRuTF50S114uHs4feYKHU32GXvyvk7k/Ja/ZBYF0j5z9ymTaUpn0wOjKM3XQ9j/YrSnGc+dYqIG7/AMS09vJ9z+TQ9AfxfyagOcYH7mcm8FfnPzLPdyt7P9mZ47UHvpCKd4vbSag7Yo+SOACdj/Y3rcMVQzKnBBBWullPsx9Tc6PcYboldj5g7HbCnzE8Wcln2hmZN7URpLfIHtEi14d/mCWV0mZAbhTDWBDMrMPSrhUCFpVRgXOvp9hzKufiV0hn0dfQCVcqJh5jpAbUDqwK6XWsl8V26/GMJw6HzM8pa4e0Nxjs8eWPVByB8MB2nl3+WFrV4uiHmqHxcdJ3A/lmZ1Vdn7lKsO2M94Lx1bKIs3SYfE1e2qiy/c3gHjH9jXgr0H5YZNNVb/LEmoXLPfSamPf8A/ssX9gYJkAnoCxemP3TALZOo92e+FT5j9if8gR1Lz/2fuXrN9NERhfYARD49nfQQfI9r5H8iHUg2eWIyLehNO3/ABkq2CQg40eN/MPqLAAD4lQgfCIC4OtRsAXtXylot0H5TUd36u0dQdoGm7FH5lcrLQPD+T7QICNAw/EEQ9ioD2hiLtc49Q+WO8dkNhVcqswu+r4g918m2gVlj6V6F8K68GhPpv5Ea+H/ABKIRt7L6fsbyslhL3qV8bR+0/Utjg+tpWVRMNC505TBy9oBi/aw5vayx5RAb2B1WjzHbSyDyJ4KPEOb2sP+ZhRvdnZV+SCjT2xDBQhoWNa7/wApdvwr/Zf+hjonImROTkIPUhL1Jk12bJ/0/wDZa/e/7CDUFujT1fLucQBEYTH0xp+r8yseAOjqZwktoEUqq2c6dzfWDfZ+Yth6f0y8IYNsDYv2dSNrwAXc65WyYZmfq948s9LET3irbl2Ida4dWeJsfqyiuE2ejKe++8PFPTzvydHExWhgDA+HuWdoWo6Mid7j0IqRCMTQvL7TXw9osFWlunTb2agIoOYNK9oOwmSN4Q/kTr5PMMvbrHu08IoIsd5kOW8MvXQy3om4B3WHwyuaNflQuC/gh8TWOTc/Pn5ikK1la+aX+Y0ryDI7mpK6/wCngjp3befcP1E6xf8AphjzFL3mJ+IhkHzWe1VHQ62LvIV8QzRoZXtY95UamDX8kPk4/NHUc0vgcfMVzR1ED30gfNd5b2mrWtB/Ipl17nT7NS3Qzdr5hVBbIoHtpBeF4z+5/JteuSvtrNQR/wBBmC8ECj5g6JOovfMWZh0X4z8RjUsYT7MyzzvKDiVKgChdlB7LBbCbYX4uL96OP7lVd7oB+pUazs8BmX0AuG2BOkG5VEq0gSruaRieo/Y3lZ9TEZjeZoBysbYrhiqD4HjO6UoH5mhe6IR4IiOZkPzGm8dVV8Szr2rl+Ie0Dg/ykQ2IdA9pWr8Gz8QLor+YRzxuEPmoPZpvf+ZsfGveqj5a7HsEdS9ZX8XNa7rPuxX7br3JMRhOubfiphLdL8QJoL96/U0zfYyxEWRsPkSUx8rp7aQoI9sHxLufk/zZiCu9un3S7byX3GZ5uxa3xNKB76PBqxXYh5f7PvOvkUOe8qgC0uV2CLZzz341e9RGB38J8P3cGmegUEWA70uV2COsptq+2zzDQC38OxoeJjv7YY1bB4RHVN2FD8fKCvXm7pZY26+2Lgl/EK8HVg258iNvP8HvKAaFRD5lHi7v7GCD693ZUOrFM9T2m15z6uOCAWDOP+pZdH66ylf7Lgct/TEFhWXQ+C8Hy7z6/wDUW33/ADAm1a2b3L7G7HhM0xuqfwbRH935l0vD9cwzNCedBpvGkeXaHsicoGkP+RHHPsEreHQYsafvakJ00uhFFA8NQQwx0CKyjrKMfxQK7fiN3o9iIGk9oFNDbs/4JXWnxMNnxKiYe0GuSqazaK7UytaPcia0/H8ljYluQnaPGaDy3+esPUl/Hsn8lr+/4lRHEwLoH7cIuTTRs+m7mziY57GbM/EAOT5IZlnHwcG5w+IikGkT5q/YbywbDfUiplDufyDbDr1r23OzJHxszeDoMPk3gh+yBUWvllhpZdT8nX2MJ7cPKNIfPSLn+WKuirLRwkGqPN6u7Xxx0gEiaBqvsv56QFj55Zgtlf8AkCoveB01TzcDIKA2U6OPemGAdaatwAvUQROiZPEWuWBV2OTzcGGkGcvQ496hR+LFImuHVE+TMTYpyHg/sYxaP8AfuoaUdEUmcF3/AHRNpreX7P5MmoNfcE/ZL1Lclid653zWsAYFuB9n8gEgBuPhz8RLmNw18ke3YtOfYahtT0b7n8gcTjb/AAZ+IoJNyz5GJk23Z8Lr4m0x0D7n8lkVjhP9+IZTPTvsxFt/Lo9rqV8qmwX7j+pbXwNU+GGGAdgR+ZZJ3eo9rqGrgNi/JOGeWfDUry9WgHy4lmJ5Ova6hSgHDPxKhFarf4NRotnBD4alO13b/MsRZofyMxphrBS+zHzllg+SPgt3T4uUgZeR+YMPPDfxBKZjptKlQD6GYJZvK1D3H7JuWgC2f5REJaJCYZlvY/MtqF2CpkHnW2EtSptAuU6pA96mjD3n2JrndCE05vmx+ZkthitHvN9A72PsTTj3oJ7jNj8zzACzYxzm9ia/uykshsc9+ZgrPSwvYjoA6b4MwzaPRPfWZ8vkV8wpM5uV9iVMc559tZipXOj31lVr55e7GyhuBO2OifyvzZi3Bc78tZXx1T7jGdY3pjC87/dTcqbjfumpC3l9zECQZtWpeNuunfQQvK269y/UcsF1Vq7rmCyqeWMyNil8nHmatG3SHXQeIxdTMoveXMuynygrTB+xBBSo+YXV0+TFA6aB7pZZkfqY4BoarXgN4ijDd1fA6uekamwKp5VllW95TBcbBQHWOdKXL6G17sd44azII53J1HvgBbe6Eizz+cPw+8eEVkeUv1oTjjacRswjtFs1dh8uCWEF5z+hwbENqE4eByXbIIPuCd4w+dnQwHSAbo3JHKKqwAWsZzAjLo+AHuwX1EIlR5RL4pdKTpZgIR+UUip/igcvhKpQjWGw/cpWv2ID/lFe74jhIWKq8l8hAqDf4ltfwltaviMJ1qCp7iaOpKjWnqkYltVeIg3e5CcM4ih35tBJa3MZ/WOo7k2fzI3Kv5IUWUo6keOTRlEpZlE3eedRBt/uQv20W6YmoKdEoDIy2MaDJ2AadmOaggF2aiSnCIQumy06js9pStM2tfVt6Oe8eOzCUfhCx7y4pSC6lWWPioPpLVaDjX7GyGWvv09zQdo0ynmWpqzlHxUectar418HxBCzpep7PkEHKmFofMJQjhFsYiTW7L7jx7VA+gcovu8+1ypFNRaHcrEbtkeVr8RrmM37dyqfJLGoaKwdtH4hRhNhb22fEwCp3Fl8cpPeIMvbBp7H7IYHQHyNHmoM5cdw5w273DMKz2RffWB0RzV9mmDuLN9hgXnHI8xZY9vwD/Zb7nv7D/YCq65A99JqB+4l3bXU/BsgUpjZ2+Rr4ljvn4c/qG2Dd5ezEOScnwGpY6QLPkqbCHIPw1EG0cf0ple7tW9xgyxFaM/2LCORn9n+xXvq33FwyTkgDLgjcWD5imBcWP3FKd6T8InS3CXzLEhe4H4jTgWKoBhjRA+YOCQ4BfxNCc1Sf2f8D/I3JB+AwtriXw7rWPaNWvzZZhTK5kQgupvxKkyu4g95o6fS79Qu25AKfEwWRyC/mCUqO176R06m+T7H9gu+jAR6yPCL7rOwo5fEpqZ3CnjWCcPwD5WLXyNP2hUUeFHxcPopoA3lZ7QBF7rLlrdCvYamPh8Ugui8PlpEK4Wl7H9lK+rB7Qwt86lzTnFQr4uXVg2c/p8RzSngHu5mT6lhPK3AVZaoj8zYrWhHdYjfVmgvfcEFcfp/OCVGsOyMll6AXsGYMVvscOQ/tIYFWaMPYY97g85YAARIEsqJUe6LUIvVa+LgoS/6S6vxB6T6CIbIRN0J4gzNUx2/fOnyYVRfm1LLMklKkWGBE9FSgfZfjjrGM3i/wqHbPWNOl99Jm+z4juPn8uh1cQrSk8rXWfx0gMDMAU/Ued+ukZqHgQOVqMIWquB3MP2NoQxqWDvpl6yj+j+R/wB5/IY0mh1uLWD50I3Q7l0BjA0DaLXHu/5ADS8/5FPePQBquJWyyVw8KOdnB3ggx7jP+ozpe9mf7YJzRt3V5MMnQAughx/OFX+ohges4AuEBF1XeX8EnE+xl2/Sxo/YmIt6gsc9Zb/s/s+x/wBmT9n+wVXVxWOZ5CZBRTZTJrs3K+x+5y/T3lQXHCf9S1QrcdYM44HVjpPp7xZ+n5mGhdP+pc3wdA1/W7MO2ttbPhLZGDmCdpy5MKqLwKiaJqJzDHr09Ntvq6PeUbSotlo2qDQCUoonaCfZwZyL+LR6S4Z+wE/ZoxW/2xwDW9MCYM8Uk6bB0Zh8vWe/J35OsGtPYxE5GZf0o7c1KbTyNYepAzqoIJxX8e6KCPUH6g6phBUcIfyJEUHUQ/kXnr0bOoU/DHCD7eBzoPFyuq2lZY8JVj3lkz8f8iQG6PhDMy1ZwniT8kFXBQUG9Dl7ygBHcT+RwpdRE9qjQJb/ADZg8VDfCv5P9LBBu9e8Fw6q+YfZLYv3iKWlvX8fsGWwANX+bI8hK9Oqpp48O6gauMg+Hb4qW+LbpT2cfMEXjkPhcPhliE+iXGLbtea/hgHCNMr7lSxTDpPth+IpUD3fsOYarOWz7yxomAP2LR/Or+wliupF9xMxdXYv+5ZhZu38MxbByfkIwo0/OX2p+Zhjrimj30l9auF/m5ZVDhAeG5Yw3DV7i/iIjsnP5v4gCW1lrezBKLsi34Mdi9AH6YHJA6i9n+x9y1U9xYNVjtr9vTQ40VZb4ovRpH4lvS8A/LFV4nb8RNnoAEdaPJg92UFa73jwRzjeDPwSmG6i+7M8F1F+CDwQcEf2ZvnS+7B3a5HfjSC0m7D8SjsJf9JW7FYfYILv6usXFr5Ss+9XGMcpp+o3SvNj3JBTd4yJ97SCtLrZU9tJUi2w0fiN9Dsp4CBrxuPhrFd2Dze5rMrz/avLmEKhObYL9R5+XQl1S+jb2dD5l569ZPGj4gICNgwRcf6qohZBdCHl+oOd+Enu8+1QNvGtVXdcsT7MrHXQbt7G8H0s2XyNb5qZk5YCk6HHvcF0DAFKljX2GEUjqD+CHZ26NDq6eFzU4Iz3abZ9d/YWqAc/6jqQqifu14LYHWYTR5e60PAGAMT5lfc/cp7mx0B3uWQHDk9+57uO8rvVbj+bPjSUH3/MqubvvmVgiuhyA2sbcpuvoS8vYdYSBAUBp+Y8aQNsP8DffRNh87REB2tDg4GwaR4U06/HKDPxRW6FJgsheDD4EPMKgBQQ7Xsm5f2RL9ZgAAZYD0MEW1B01LuRX+RFsUeCNP6T+RjICAtBjjrEKpZRoAcQzfo/kC/w/k6yeIlRveMH9Qpx7pBdryfyf8N/Ipn4f5EHJMbh1jQQ8SzY9v5MB+Q/kd73j+QAuL/IXZ0ejESUq3LqbzD/AHpbf344asYeoE5Ha4teSCLbcQMvbphdYROQ05QkMu5uq6P7D3Qk8FiYJGlZezlVC4d7ymsLGehp0H4hjqbP4V9x4uAA2ecApfu4jYLEWkpRarS3lb6+yCQqYVXVZQ7Z6TCZ+tv7Aulvf/YGBWQtcjdj1IjoHcgfRXuhkD298Z1OpZBd33/2Yt/dEarceRNezcswAb4bravCu0rx7kW8KyQmKtVOQSVbVvOe7x7VFdAW++asPFxRS8BROEcnmAv9TClaOSdnUmpcNPbxunuxeADX9dh7QfykTXeWZpTMyr1DzZGnnGkAfbUZg6PaP0HkIMSdwYiU8ICPiPDNvW86H2izGdk90x8EMPlifMHvUwUzVET01oTPvNvIe0SpS/TqfiCac5/GWS/FdJmY6AAPOsfdyHyZ+Y+TX4px8wwhnjPcxLw53AR9bN6/uSq2OMffD8w0juE+z/ZRI8aj30+Z2aMgjnPUT8Y+xU/Ipm10+sagLsDLcPfSfOCiP+PD7adz17T3ev2MGK3S2/xULwN2K/gg5Debt96hYdeK+1TUfqU/MvQqMl376TIOnkD2JWOyWRnQeBL7Rr123E/2M6Syhfd/kQ6gB8NJSgBsWQwH5i+wgjzkn21iDtzfLMgdel7sdpSdmWquMp4IJzvl+DMWKjbT8LfzK1deFfliDk/L+w696NXwSq6PH2B/MWttvXtH83PEwI+GYABBgt/YFNbRD+CZNumH4MaPLBLj26HbQe0AAMNAx/MUfX+ZUYbSzeDTzAg+wD+SnzKCE1tXlceI/Y/uNdft7zNgbr+Bx3YCqHQiz2Tx7xyLcmnVW2dB994mJMFtDy93YOrUxre2Y0cavYUd5SNNAg8So/jE/wDGVqZgnuWnUY6IqJbtZv6vtAgQGwZR/JBH6kfkmwFHm+R8Qc5qXAPsnXVhbp+D+R/xz+RD+J/I7YFsHKSsD50JgMxZ8LA2Nofww/kf+R/J/wAF/I1+jSEHiaBpy1CnlaqV5RWVcsr/AMf5Nz8H8lH9z+Qe62I3y0xZXlABbeAAKDSL/i/kD/k/kf5B/IRhojcvySMAHvS8A4sICQEsupfyBS6/OB/3ygfvxP8ApmYxnat++aeYB/YwP+2P+llDRO+CLrMexboMutQ3V+cLV7+EKpNc405JlklC9UJUrqdT2e8tbWobUnJM37cbx8v+xTDkoDqN6xXfLj+g+TsgG4C9A7jcHXa8ojm+7+wqj0lSLNDZbDdNx9zrBnBdmR/6WDKOkaveX8NxTK5HUepEbH72w6Ozpr3lCQaGF5GR6MK5KaSG6MLL5DJ4j7CCHo6edPeEisVabhMkCNTtiUNB7Sjf4YQZjto0rB0/IrvFbKjQXw6nUsgf85aFH4QEJ/pwZgVkNkLsSnyHeMaJgLd9CmIMZehLav25TTsiU+SOaf21PQq9yXsHVJfY37qgU3WIIkrKT4S+DjFJ8kHlK231dRgimGovzh5CHUnYJGurDxL7/wCvEqani++Cn3uDa3Q58OHtCFe0QKdzUlbUOLIjTP8AqibYGgPgp/M9zgR7YfiNjTVK/DmUqXHqRHlH50QFrmxB98M26tsvwfuHgvt3+Zcg3cCMsw5yPuQNaHUB/fmPlmofZ/sHI2NA99PmWYLoMdVyDb3J/wBV/YQSVkJbn0huo65RwupmHuxOjm1/iCW7+sFBC96Dn8RsAcxRRr2+6VAiqdby8BXzFd/eKgiiuqLP4h1gcv8AmAIZ7r+BLCp2UvYP3NfzX4oX8xhXXhy+agF/N/ktczfewEDwBhR8C5lvXVnw5feBR1VZe7UwaHl/IDazos3sVmBZnbrwFW+00C5p9/V9yXIx1bW92rYozXvYuN96YY5DkfdS3wMHUBxZ2HU/EPk2o293eIf+4kAMq3iJNl4UnVwRtOGbi+6y+KlkO1stcrq+Yg/g/wBinX339lcaaM8+aHVqVk91vFxseHmOwysGpyt2veU/1/2OJfv/AOwAzaURwDbGoekLy65S3l7RuUydL5Rte8pP3P7Gn9j+wSDXQB8xNIlimvrun+Axi7Fs55G1nSfrrMF/f5lgjPvmZiOrchl49DeWCV3iyv2NDaIGPs7w3B9d4lqPvvEkEvu8mw+dCKr1zegOBoEp/wA5bNP/ADiF3Da7At1YKcxQEL2Bvy3B9EeM6/2zqvbGRAtBgj/jLRhcjyPYIUYDwn/DfyH3z8SnpfTiVg0AMLztwJx+3/E5LO38TL93xGj6viJBA1UxS4jB+Y/kt/sfyUb3k/kxfofyYwsptupt0TzFAQ9aLMmku/yfyX+j9RW/2dokWrwtbJjUafE3H+vaugrzcCtUovdKjTXKD8EEMmdsDsygVrVPPybtzEpTS3N0oaRIT96Cl2V2NdohDFQ847nPtiQrZSMyX86Gi2v01lApI2f9IsZFSJ0HsPNzTbbbrGa4BA9/q6wvwv6czGIp9t4MJUiRpoG66TGyzCy+2Ta6OOsDWkECD8wB9j3mt9jzBQOrsih+HEfo3xzrcO+j0iXDB0JwmR7w6zyj1/lhsYbWtcjqPUmTEd0g41fY94hNFB12X8l9IIIxyeiEhfYo+GOXg3Rb0s2eRKgADVncafA94MSt6NdOkq/hFyhhEIy71FtE7sV7Q0ocVneVl4SDmj+LvXxcKhQdkAHX5s2lrk6Yj2I5pfZFOgflQccqq+eryEJJWlA9yWGPbTPbUrB2TJNeQ23utfKHVHE/CfZYXvX+FowJj2CdASGxyV9vygPacXelv5H4ilJdX8wh/mAn8QpRtQEhXP8ARfxMfERdMGv4PxM62G+D2w/E48ah9qkr6K+kvT7uJmaJXAfJn59EHDbFgvxMylzk+8qWmdYoDlu/iJOxi9i2WsG/9htgh6Hr+YEAIiuKewjgm7PmNR00m3zTiMTl9We2kpKWwkHIJyhNi1fhxLyXrCivg/mGVzlXtj+5QE9AlLd/t/YI8pIP3D9X0EJ1Fcnaa93sB7pv2qPdWUr5W5Qfy/sEtM5U/seadVj85o8xd6iFJ70fMMgWx8RoeCYwduyY3X7P7HZC1SfuWtjaBUchr7CErDugLwc+VmlCQAE/5mBZftnQ527hoO7FN2OmTONbxTvD+69Fryuq95T/AJz7zCFBsUCawtpLI51HvQ7xkHcZ2js6FRBwJavt+IDU/vpAGKtkOgod4lsrcdtGX0IEBXx/zKfq/Ex/X8R7oKkA6tQOkzQPxy351doAO8KA9pj+v4j/ALP+TNn3P8gSdaHyMWB87ReEWj0BjA2Jx++/kw/vfyc/vv5FBJUAAarLMoE0tFHXTozAmD3Mo091hT+1if8AVigC4N3fht7wEumvAFTD/qHD84Hd4eYFK+1mc6xrydK6XcxP0v8AYPA939l3/e/sbn7n9gqyY7lZzFQ/N/svZ9PeL9X9xs+/5jqICOs94x5GX3fXSlPED6P7jT7fzM/p/MUv7feF+30lc6srz2uFIFeREsdYOQzcQVLF8wCxWuK1t5SxeoRdg7I5GWb6DaDft3PMH2TQ0+2Wb/DEmbm5WI5SsDk4+nRgpsAJBahqJuRou3smWrd6QbCj2RGHYB3I/rRj1jAq3oH+TGxAsaUkFQ1MDT+TL+cD+QbTcEEdqSUlLLO38i6ZI5BtnD12DqRfIvg/kY7Osyh8RXVJfb+Ta0NL0QZOjZF6q5rAOx7vZBm/gNnCVY9GH+C/kLNTw/kYLBUk8JKhRrsP0P0NdIjr2gWnQmPZA5pZaHzMtwCs/EM68krypV7p+Vy3jjmqfTiH9FMvhvD4uAcq84rU3vijfvA+YoH6G+8WeEiuhmqfNeHi4VhmFe6WSDFiecsZMeqOF0/baz5ho1c/h/cS9ajV38tXmpVqmix+Y5M+/ELz0UwmvKPeoT2qGkTuPmD5gCL3Tfa6PhgmcaNhBiyjlYjSCr33wYKvYlT74fll6g3vyyn8w70HNnZqUAN2G5fT+UfMWp2Vwe7HxA/Qf0h2l1pDUvxZ+J9z/UuAAJkD3Ya523+Ajlv/AHUYlSa2ISkbEe77LPBmBgAtFp7a/E147wfk2zqgo+Rjt1CForvE22K/gJRyjmex+2DrF9sP3KipsQlrRYdYgFMrREHQzHF6vHzMoR/0mDwS1hq/u2niBf2iB+6Nw/cyUF99F8wOXtFxDc4z4G3yw8YcIT/jpwvwleIamXeAZZ5pAMdC0eXxAFN2THoaeBKv4oZvwIL+CWgLShnXQHdnYrQRxrvaneADbahbyuq94/56a8z8YZVAEVnmTjrvdLTObIVH9ry2yoxg6JRf5Y/6cHn+apFqg1Tl1NLyzwS9LLavMGV3iOsHiTpZem52bILKzPqalvH+C0OsHCgCsL+Q1he6a2Xugi/kTRLCtob8R+dIswxp0BwNAlLr7/8AJg19/wDk+n+Uxl/Z0j01WKtYp5OkLUo+AFAYgu33dINt93Sfdv1HCiGfsS6By3CDjxvh4hQfa8QM+17RSE0/swsK3X2TDYyHbK37RP8Aqn/WxzflwQ4O6gGg26ysD9wkGcvXKQI/3Ru4jba2S4OyxuR7pZBJBeAf+MaMe2f2Nt6KKDhNZhukXM5vera7VBbr2z+wY/j/AGWXr+P7FIVXy/1DMoNQGjrk5N4XhgSA2y5X+St3u/8AUtrrq7v+oDdCxH+p/Tp/Y1k5EBc57PumNEZNxBfzvEjC/TmU5PudYKU1/TeZ/qVQHZzNdqgw8o5Orwwk4m2DeIyJww780tGo5kMuXtlyO2NyQZGBpoVQh0tJyZ6TZXM2uibPRlmDvU/kaPs+IQtDff8AqLysxe+yqPRGBIi1mw5oU6tjtNLbFZ+Jn+/4idrv/maY3NgTtUNg7bePVFHejKI4GR3VHuidZtIdVfBD/R/yBvL1/wAl0j/RiCDFvB0H8C9osjTru6oX5B3mgmSsfJE7ImuUpFHuZVOhDZ2hSe8LgNto8DDzcFUA1V+UPAitHpWfEN17GWzZ7WNP7TmrPm5aUrV/pcxi2jW/5qvIRzatGp8MLarez/YpB+pYMumJ1586ntFSjbPR3LF8ELAkap9+T3qAVzoPhgpvd/8AYjZdab5Ze7rn51+Er0OZHfyKfBDFp9X8gfmozLmtR/cDJdw1r5n2/wDYJm6pt64kRjVWOeoP8zErNh3vgf2c0dfxJn5nUDA2+Yu5p7S3GINbB/bmJUyf/hmPmCj5u34VTpDMxT/CCKBykcUvGTHqmDyw1xNx8Zg+YEGejUO2h7QSJaAAgXPskOURWtEuFaDje+g8s1cOyQ7sPAy96Gcp5dPEOm9kr5+yIsidiGCWp38DyY6+XAp1CjweYZqDcs8plm18Uf8AMje/FFegtT8EO7FFZeEpxrvakFH2hS+ry9Wco9ons9oPZ7RuzaCdQ9D1YGuuRw/J24OjDdnQAdAmLQnAPaE2JQe2FwPA72eCU0lRS7f0DioIoIBijVSgziorImTo5trliSijCkeMddWMYJdRTWa5Ase77Hdh2dw/K24nYhV5gEogMQ/3c41fQyst+czeUT8HBKO0RAK1jW0Q2jA1MfsW+Ia2O3fcXVbZRpcNqlQ1UcWnOaqX4XBioEHQExAJXFRATHAvUdCwz9PfghiVcQmI7x3tWrTzYhxOwRLhRUaSUHWIzUGUXkxjrdBZ7TFQyup4TqNkuyYWBauULzRdzMuLYi3MKUcx0IyjHumvhi4rQIJqj8O8Cm0EHSWc+hRPZR2DuddSPGxHeQ3NkgnSJsSojSyL4qEtKb4fZuupzASOjYD7vtqSvqVFLIPMs1AQ+PkuMYWQ30NLu16xqJ3VjpuvHuYXACxGDzzE5hFdRM86qB9FyX1lQJDQLXz/AHTrAJRRUSFu0dZoc3eOit3Y6iLS3/Zsmi2qKJyjnye0aHRrCfhMj0SChi8x/wB2X6+/HwPLanQfAY+0M1QDqn2E7RGTTX947kx7a+jMuOHwjTUOyIGE5530eQwdZrfKfceQmAOwQjoqveHX7IijB/4Ji/Uixv8AuYi/NxcD3HV0w+8USy6xXecPNTrUoGG4vCUMh4RmdS194F8zQ66G/CfcY6XmpPbKEKA7L0feyRJ+FloZ/MszbMf4U/MTqA1DPcx8p9q/cPVROmvmkojI/vfsFSpgbUn4mr6PiVKbWmfiMU22ZD2VHJJ3HhwEYseu/AVK890KD8S/T3P8jpi7/wCRE3MPYhAxRVrR2vywAPVonxA97gER0VD4Jx9//CNp97xBiw6WF2AtlRVmPbtbfiO5rW9Pwy+VmlGAqD2I8j3sXj72DXi1gCJLYq6j5mfFxRvawUOFr8CEROjAiJoRh/XA109yKQhiqedXkzGTNCLiy06FQdxUB75z3n/Uf2f9T/ZuD8/7MIkGGcA2zPNGL3CBrtLZVnWIanKW16s1fzYdX5Ef6xBSIuhCK3MocPlHB5Z4lDArJyQbXvKq+v3jT9fzMmgffMJVKvreZecE84N+M03iA1J7qC9OAwQ5Dw/seF7P7Oj9v9lBv4f7NW0i7Xew7sp2oWNDg2eJh1+yV5v7JefozBCZsVtTgMasoPhrq2FVjUZTX2PEWMex/ER/j/EC1Hx/EoXRXT+JYaNBQWDGxRKB+r+Ti+P+Qbi7n8lX9j+Sm/kP5GtVYo0V3pyzXk8P5Cr9b+T/AIL+QY59p/Is+78SwCrRwaR4jKWJ9mDjLTgN2yC63eVSgLeJUP4ZaFmwOzEn78x6nlFf6Jdr7yFJKROtSrXReNfeayaDrEbf9prUv25g+v0usSGX6cxCvPUlqOdBowsU5VK1C8I4qGf7/eJ2+vrD7F+Yt+n7wwmbVPw25NyNQjvELfv31Er4Tz/sKtzqv7C2rvl/YGavd/sQCtsVNkrUepKyi0Ij4J7DzKDiWkORGHDfLKWy7zLt33hj1qwPDL/Tt6+/l9GztCGNA3r+DqKR1N3iG57EDuvZgCLDikR9Ae4dyYe5T1hNrfIPu8sdYSybEIOiQD+WUMe0mj+BKBGWW/yD93HbH7AX14YxwT98jXuWQNZd2I7h8IGbvZHyrY1OzqQfsA8b/qRYrxgTwMeBFiKsqR8kP85DpfZG2PyFEihHmzN62ewJ7FAo6tT48JeweFZ+Avxc0pjtBrRO0UKv8RPUmbfnaX5laP8A82H5JRZBT+0q8hDPHiHxBGj2jb+iB5c0LTtqI5AJp7Bse8wJvar3xPss4Yax7QMTQDpK6Igz/wDVFB7qkETUf0IHtNyLUPlcHtBlbuv9poe0CxC0MIaq35nWrzHQJ6ZvsMwHK+ie8P5VGx3d3fANvlnQ2oFyl6kTyQ6jLUoIJS4oxer/AKgx1KzU6/qJSpuvd3WY8gRBqLygzfJbfgMr2mQG22iORz7iDSWRcnQw829YEADABQQN0CusMVQOWX95VGzrfkvpE25ZsVcfiKJp4uMEomsS1qFDmayqTGeDl6EP63yz6d/ZAQd8wlodCiFEazOURGt4lf8AVoKG2g73sxvE09L1PoVUJgo7SiakDmIws9471QgByssKCjs25uXydpQCc1Hfq9YLvKVr8xBvAOpHMpWMrm2d2IgEvQDYdnjfWZREDaD5ieHvELw94GqQa2y0a4H6D87KEAGmYVkV3jcPcn/SmQwd4ywoetwfyvxFwRYOcpvKzS/NFP7Jq6fMdz20tjR2Szg4TVlvxB/ww/wMAFdth/Zz+y/sAc3MqACCStd4hBwBESnPSC1+x1lI/U8x1wcf7QE+97yp4PszN4rVqxpxZiAsLn/aYvu+8GLpfXWH3N94iN/R6wkO1a3kM7MRMLRDAC3kdYkYAurf5lxOLMh+ZYIT67wNVBx/WK5V9f6wawh4bio68DUmG56R/ufT/wCZz/e6wOyOU/3BDccn95gEFsfS1hlaLuXsmnuOs6JFhntE3YeMuTKdEbDDdKvmXsE0uv5nULikCr/SxYUaLug3r3MMQ6vXDXa4Ia3jOePZAyi9pdZVg5I8kTMVx6NJQ/4QrGgEpeMk1HQnTviWNS4FxRc4kft0zejsw95KCz2HejDIJYEecgeiHmVFkwtC6svLxKlI0ix4aivcOkgXgkOqIS6+RsXaOOSVKTgvxveP1eE6u6DMFoycOQbJD50JY8kDWQ7yKWuKi+N5rW2tR3f4XHzZwhOfmE9oga3aZmi13IhLgyutQjoxt39pihfbIObTHiUf1auLjPweEaMDHiGDsZ7xFl2rxCgraRt1Ls8zKJNZE73FNhwKLvWkM6q8+YAqjhuluHupp7gIA9Ec+0v75Qlr3z4hdcaxJ4bSnvCeSABGLjDsD5Y5/KBS7po9vSVhwdbTUtcoUS9ujR/XwSgTz86Gr9o8H8qQPmI+0nq8NOI4vlHYMKRfxCk+mdx7waLbe1NlvaDAKyG63X2peEzMS9Fph1KsOPKxVgwKX1Ey8Gqi9p+WDlNExzYNXHQ6vhgkQ0p3RFvNQzrhQhemIGpbCj3IhuLZZeoIl/ZVzo6PlGCrSsBANxlF84svAxNSll4PqFAUVo3zzn/5R30DXNM9Cx76Y+UmterRZrVPYKm9ON7o04jSIUrvFp5YXZTBBzQdnLHWd+FLyOQNODXK7JsTcqAPdvpDVhnjBZK6wqMV3yA1HrUGeAtVtgxdWZTaF/toL6BLy2Y23N/NxkMSBdAg6EHZbD2aYgdBZrrCdl8iWqslm6ipxssMI9izGC2HcgwsQBJcA3CG8FKG63uu/wBBMCEBbZ0Yq4OLKBWHa5kxT+J4XB0mKiII4I+5md9/+sYvXs1Q/LaXNC5WMBWBUQnpnKctpVgiwFCpN2N95joE0FsAYIHfuR6vRS1tO03mrI9RZrLvpNAUgR4JoanecKCNOdcVrr2Jd1scIyvUwILXvMfHbNo9ewQIlS7ClAZ0MvOIdaJG5SxA5W/1pOdgvmOYgq3+sQNt3/pLRR+AF7nSHmPgpgLdcPvAVa+f9iz93+x70aSiTeeAlWt0BaY5O/6aiDb2hZG3tRsD4gjHsoGz6zpDiJTqMENP6QpdH14mnpPrpH9BAHSLW/KMsYYDqrTZPmYpTv8AxiCi/XaOX9UvYCzGb9kb9b7QRg/rxKmDB1OyaX+SZtDn24brKXUXsfXiJQsYdiU5qX9fhNGyOx7MJJUl2fxl4+D/ABg4qEN3Q2L9on7aMhb6aNyJ2vvxMMKxjhEMJK15xFtuVBNbaQHJiEM5QhONJrTMqt31ujaNIo8OP6Jwd6D+RC3yRtwNGBoMIS2KtOsEVZ4B3GJrIGoQyjGgO9vil0vlLwh/ygs6sAROSGvCIoFkimGm223EOSA63DjXRNnowd+0SH+d4/zqzrkMCFwysy3Qf8QI0XTRORhGbq+O1DU6M0F9KHI/MI8CmRTcag94iW8x6h1PEP2t8faHZ7o2NrIjnp3LIKN7CQ7kIHK7TbWmB0bgP7xqflQt5zVcLkYjr6l5MMniEpbbUs40Hwhgm2wHrTh8PiH10twnfUS1EeUTfk83MFHWmTs+UIrbOavU48GYGXgviMnhgIgze6AdTyMFuUHvI1p8doYFjIQ91mIU7Pz7R5DGyqugdgZPBMCtMiv0KYmrcxE7w5+Y/wD9b3TXqeRhjC5LDy1p5CanQlpeKdZr+wI+EvzAgI6YRxRnyTuFvzyPeoS0RFD2OT3jahtik6ZyHvKnQCRy6/iEa1hMXjM+gfuNuK70tuLwEE6NZW8FkFV4RovIMpk08q19KMp5ioUZInqrLEBI1hDu8R6ljp3Hfg8E0E2X5i6eI7p+C4PAIi9LQOTUxGrd2D6Yy/EXEDKKerqfMrFnAO+l7wxwNuJwvB4IrGja534PENki8x9jWIj7hd0Xr8y1Z8v0l6vioaVsgi9V1fMV2PRkXWseVRGu5QIdfwLg1sx3kLMY1tZ8QasDMF8i1fkfEQqMkD01XsUQ9m0DHnmGhuAqvgcsUWm3xjcNPLMH3dLXK/wVBjbYQHdhQ7rUO+onVogY3CRwWB0gwg4oX1Xd7wWD7BXAar2ghcVeX1oTRRR1TcLlPwRMKtWld0HsDgthVU9oxNIm9OFWnQ1g/wC6KV9V3erK13EA5WKweoA7h3S2HPTyWXQ6ShE0gWrpF+SPngNDprHdxwDvsWywMoYHK5N3rB9sQxmCc7hXk+I6/dOzqW0haANf3jGbOKFEx2dZqsJQXtB1Xywy1Xhd0m6wBip1jIQcXPwSpHNSxc3fmIE76lsvu1Dobo81iCa3GvPau0F1uZqrELauHQ0Iq5D2hNr+bK6HdilohePXF/gg9VsMo8xrbaVlUFmC2ozdcyAuA5zjxEWdSRe6+DEPI/JsIAgxwAXBfADyp0PEbC+TIkZf+etL/wBNVRNLEsS0zaiGGFmit2bmeAV+5cy+RGMAoRxqfuY9VamR92pQewSj+2tCxhAO2kpRmGVFaAvMCLrYe1IJSOh+EZjuI3Vh8LBKEAgFJPFXq9iPLNWXINgKluQlXdgXshKuRsYuTAkphRuB9lhmxjmQ3j2lamNBwvlnzGK4QJ/MSShDl6JRyOYGTplVqJTTSbTChG3Rog04Z28q7/CALE0CtG70dGXrKlKJoR3SA0Stt+40w0eg6mDBZ4WldKctt+ItJVCtIDvI34giv9x+4p8ypJJArYXkTmYHIIIXivQP+SvcC9B+YQvOL1ulBhVnZvVYym4XBjVjhNE4gfLjjaS6S01Y1mKYUFTccEyhO3Bzkuukp8a1x3FMQck77Vo8GlvT8AM8kuCCgA+ULR0cRwn9ELVCidHSCiWTJ8gCTWh2OwerPMwIvSsY2aSpFvQN+xbKCiyxbUwE6OIqgS69oldpbBXkrhMQUiS0o6IyPci/V0ZfZQSiMUA91R4qNS57VN2FpdSkr3j4lscdGqzuDL6Qi+qrZXwJCXKpKa1Di9gSqnm1PK4IXYoi3UB8LEVH6Rc4r8SrJdCeEw8MVWRal6fICCa2Xk+1NeXvMHQ1oWraNcYm/wAd4QIPaJU821PwJ9xIbewdQoBZfUjUWVTh2MotgtkvyVT2ioFDuIryrvHfCCn1gBazyE2GOIvsHzBq0X7OmLwlX3gUfBeFiiUWNbiEV5RgtnNlvIxg1udGGKQ1N64V+T3lQyaIybDITTMpi5cjdcnyMR8UQjpaeSWmGNS8AFbysElj94ZT/j4MO4VcviiD5I50bFHr+Sm1twVd8Z5IJsQGuO7YmG2YMPHggAD2miS4XOmXUSx7w1lNKD5gn0WQ/K/mfwLuqUpQDAf2wj7yq15key2T4EdAmsp7gHzc1RuKeghEJCVNPcgntcKuqKAOyHuYmVF1mXlpyyoCwVuhBosHRf8AZGDVOuM7Rqb7NTj4MqNQJfMQpa+3oofYQWM8+SwTl1Y+yweZ73jsUTIxdSPNlPiaVMM/0MVe0RrXCyGjatdWpZ1IYPQmeKlDoKiRwYEGAKlvDYofYgLy4TK2MPdl2olKe7YwkQjOCHiCukzuqEB2LYZJb7fQqL0TEkvbe8sHgOhYsnxCqeQUxw1op0hlJ15YtLuEVwOL8UQubgtvFaoASxaTshfdHEDmwQEhpuB7JjrBbjC4yl3LLyxjBaXW3UD+XM7a8370YjdVCHhRBnCDGgSgeiMd0A126pb5m/plK8jT4jzldytmt7sMrjMi9oaKRawJ7UNDSZI9S/y0lJxyE7RWtWLJmlVo0C8HaqmeSNyPZp8SyZCnHRq7ZfyCDcNCNcvmG5gQyrBvY0ieTXLm96llI+uCcKIG8Z1P+xfUgcBoVQ+IZMmFN7kuOKSOzs1aVr7RKOpVYmg85t8SlNNh/KKkXYv3pHlCEk9GwmuOkpsDnmuAQgF6fNLMdrd0gAvaZOIrtW0GxmWpp15WM9ggdXf1Ei7JFP7ER4kDZFJtu0y7xwphkbXvaVI5t+MI10RrCt9OkoWk16gpKgtAdQmNKs1BPuE0YDN7BhaddNoE1sNYi928G8JEPiAqljhHRgpKB1VjhXiXTt7Fu/4qeJSO135Eem8iDPaptClVbN40z4YUb4YOntM0AOKmutqjPyeCzqR1sMF6nJ3WZVaGqJGGEpe839RR6q77t1EHW1oHeVGpDsAcBGh+NsTUSWGpJ382m3KN+zhqhuO/DKIdpQ/lGTypKcgLGJMxrmXaawWAssqVXiWGhAoHaBdw88iLHbqLNzXqfJB4wy8nPIjIS4S49yHhFnnGCuwmJcAuhdKNzqRIhmBoFg4SGHkJwmuez0l1mxOPN6PmG626YejAWLabwgH5xBTloQewT4QJY3dHtApwRKDKoDrjKUXpouNhNDDMEfl+jtDCj5kHrm5kmcj+hqnkxnSI+jWQvPwmsKspEsSC4AKRNZlklFPkHipWUNk8j8uJjdwuWcC4/LpN7ExZ6H8NkvFdcDqX4GZzCEncLzEJiN6iaD3jUREwbjR4Gvk8x68ZBDkNnyiXDAToU48Ig3Fv8zS8iMIg3qVc/wBY6wQsapNdE2itAiZHIwPi2lNvKBT5Iot9WE8WsfEpuOG4XX+Cw9gcu3lo90XaDMAcGJeyPmrRbXQy95nikLYkwdEQN4SLyLRSnq2vapc2gA7H3HuiOjal2+5+ZfMbAfgHivTYp21YnnkNUl+OMpq/b5Zow4M7xjeFEws9fIjMLvxu8HSjn4h1saK3dq2EFoDljpwljfPWDzKlhxS38IswWlzOpo8IixeSzov+DA6NCWx2qX8kLI1lKPS9e9wCjUMAdCBLq0gHvFJZaeUvXxcOomqp9F+SaARsDjg1YOjPhL0c+8XD5cycYVFJa4HnL9QOJrtQIE05rWfTOCWHjZgN8Z+YVgiq30gZZlyGiEDjogGs73perVgssoYDtKRj8fYB0w0OriZEOGAXoOgwA+9gvJ3XqwvSDctu3RBYDgU/VuzDEMYhR6NiAFQQ27whWmLQbujfumC3Z/ECOusSwK0hQ5SC22YZjrWr0jKAvb7Bz0JXjenm5X9SlVGZgToHLEq7Ejk/tD0foau6bryxiW0Qst02Jd6Ftb5LxywsVFvA14uUHUoVQGxMBLxhy+DlYkkVD4Hl2lXKB1lsQZFT1RsEtKwLWnVBztCLpsYuko2W0AMyghLmBli9lx6Ne8uQ29NI7AN1REcvZErFY6oeZfCnrF0B2/UWr9hDSVaUYrvC8SnecOZGl6B8D7wCABQcRDqgADywHXU7FQq0WbLlwmP4Q9o54rCCgM6iUdKlKuWE2VsbDIrBZDUIjclWJ0uy+lwo7K8mB0zoy19ver2GFhY3NUiMOtYgNNUh2BvwSIrWpQC9Rj5hrpKq57LrtxEBPtagGE33PMD7sJ+EYCsQPDHUIaC6Xf3RYUFdHU08aRQ4qKNEqEXxvAJdL1PCwwu/WP4zu2heo4UO8x6EXJHSqF+JeGmbUiR0wYDIunQoK0IDYjokdLYpk50XhN7NqnSjqql2GGlk3F4iFp95jbFmIDpSlPhh7RwJXsmyTcNCEbJsmICII5s3h1aldYzVZEdQTPjeWUGlQ9gDValQ9HUQCWvX0hYLFx+nMJItkI4p1OJpvjgCeE9IXyQwqA6wxTVgTsNiOkbnpoLdRhWuly3l98G3XVvaESREpclA8sZwN87hoNTkjAD7Tv0D2mWIMoAN2LA1vYmay+JRxy5Fj7R9hi7AajrbiE2CyPUfKYlcEYEi+WztCgJyjTdOD1JRKh6yisNV1let0IPobxA2IVijkqF4cREClFSMG+P5mWBoozkewdSU1hkbjgdfcuCTkyo+HXxHiMNpGUfOWyshGcdzrMVbUMegqx8Rf9AxMYCKbeYLXKsi9V29lS6SRoDPAfCNHkyB9h17ly0ykVIxKaB3dJYZS530bwsJYZ5sCH5j1AYADFE1nmpl71Kk9Wr9vMu0TF8XgPJDvC1PiNXi4O6I6uGcAdl0hpwZa/xAdvRYyJYFaI0AAqjNS1tMgo9mR3GajNtDpaqDqU1Q9oqRbRxbD1ME0tVV12Ze0skumh5E8oRPy4eHWx5xAsJQULXYDGlsr2qClOw/SWpq6LeBBPaA6A6jfscy8a7q+cvErAQaqO4pfNSxMKZAdcflH1xjK6aj3O0oNoUClC7HmWIaaIXwQDoR0zRD140J5l6hmv4xfCgSxYUxfFgj4YkdJVx0yHuhF5UodRvcB3bgnAsgL7ls8IlWTPy0hOaXaDJudydgYHaEGC8BL1FfZJtr7l/cHySorUAk94MOoQlBqGp1WOIONHf/AEXvVI8yCmsLRNrxGDJjcN01L2TWgk4zejY+esHVy6gvWt7VFDQ9mfksfBFGK5CP0ZCEnW8I7uThVYvo1Ya7KwrysMKg0qtjG+FRmDSzOmt8VzrHRBwhO4G676xvs6ue/m9/CWcK+jyAzrYs+R9yEqUBoNgHYWZLyKB2UPlgxPXIPSrHdY/RPkBo2rOxawfpWkHWy88sQ6m3G+yp8kzAjQK+d8MsNeQA5oDB0Pp0VlBYcFwauKPBtlo9mMtYoEP+ZTBdMUC3HQZWhZTDCslvOHdjLdF7b3rAZSDT9qn5GL1rYwGr+FbMKHu/lq0t1cDEeS7yrxB7puZTLb218IN93Iu0gzkrxM6wushMPgz7TdUNH4BjnntBJBrmRaha0JtzKPYcF0CwrjghksNbX08CEjNu6XzTh4Jf6NgVqOmiizGW4AXenTadoUSn5Eciu0/In4SN5si1Avo+Y2hDMNVACuvxCqodRL532CFArOUvJDwRSFCYJYdEYwXt4A2Zt8RkGCVRlXwwgvfPaoEgi+dST4I7jYwYJgXRCJS46j9x8FQutQvbe96gl7Mg0zU9o7QviUOMjrze0fVSJ0wOvv5iSrdl/O+ERDUYiVVtfEMWdUmcMc1awfQIWT4b+UoVamxe4/MNQwrhhoNYkSzQzuYepLJXkB2Z3/CLk+On6dIv5oJvjOU9ajZqa+dUWWJpcJojrU305nOyLF5W/MUMipCxOJiSu7n2a2dojuYCHonlEYoj0BMOVPkhD2ywGgvCcx6ZLcC8BJ2zpCACmbX7LXdYRarUtu6yxCKE0R0limtmjc9XpvHryhnFzQ4MNZApWNrT3g6S72hhoets5PMJbF0t3+YWqDSR4oE73K03pJ8yoRzT2Y4A3Ousrq+wJzWFJ0j32O64KPhxOk9DOlAEABVDujfR7/MVYURPg0B2SH+Cy/CYJicUh2f6MYcymz8q7ktNTQIHTZs8J2mdIFR9KvYpKHC3kFbEW+8J9OLFG2EPaCNpRj4hUpmxajjuceIMH3bUvGh7+8EKcLqy9gt43JbiSJHUr46CSo3oVQ4buu7XaP0K3Ca5PgQ2BaEA9oK0hVPoVDqMcnmiLfyx4hwKqrj8nyCITRaL3hDxBtCFuV5B3ydoxiAu9cixfiU6K4AqulSnSITYCixmQKYlDzRh9opzIjBnGhBAKtdth/oTqePGSDU7kdg4X4fXLUqCfAkPbSUcxqzAezvnOo6xYt0exwBBTMqt9YH7mlWDPg+AZhSLGooYttfyhGJlkXs2vxBer6sPLUoVDtLf+QBUXQV21SzEnAORZZcj6Fy32ey3iFUWccB3esK3OG2HQGjzcNSmUhnu6eIHo286RH/IPsbGD3l75oR610MTjtZm5C7oyux3nAiFJzuiIkOIQG7RsRRg5SbO6nluDAACgDBGcfEAu2g3dJkLw+Q0AS+hpigdNxNOW02bs29cDTuyjaYp5yrT4mkqJV+2T2GIe96DQOhFRR6aGFpbm11oRdl6iIOi71uyrIa2hIevTbdf57zLfN23cKZ76TOgBM8w1WUECeaFJVydEG7LTl+ZeJgfKqwNgjO1U5L8B+Yd3ZPTYNggAaI7A9P3d4Qi6xviEqAasovLjLDt32PMKFMOgD8vWC4ALVwBGfHisfptEwHkGNns5hkAAUAUBB1aSgm8RZo6BqLoaviH5CGmd47ssJQgsLcU+A+ajFLTGqrjfmAc64OZ9sHiFTEwlAMJGmtT2PvBv2jyj+VExxCDCK5SqinTrcNBgz5rKHbZ5gveo6az/mrOFQYmdRhDUhdCuqXfoPMsRKsMH1zUFNsv3LKjfrCLHcVn96phIBUNRyOJehyTajY2bn7iFoNDwwTuU+I4sfMqJMSMBqxrffCBxRZ1NPGkYcOkIwSAW6/cNTqSh0iFFP4kAcCLu4oVm8wRSuliZz+TrLFcKqMFfz1gv+zTER+cuwMYOFQO9PJLMT3ddnq+I9UBaHHZzB05QK2KbfuP8T4LJz3hJBHNmfQSWYYbzraK6PDq95o3w9yCXSTsehQy8zpqSn0Sq2un7ia1RS69D3ozW5MM5NBuBqMMsojAcho5XK1HqR+dLZr98Op7SnB6GkaY57PxE9ijpromzGeFW5MOlhqYeLl+u/lS4RhkjTn0GpEDOuz7b31jtpRQPDhrbDLwvpXYRvT5IFfWUIOcwG2xhYllYFVsR07kzgacz0JtCr69Ymm81t/jp1OHtBreil7X8+8bB5w2MHPI5iLC1Avba0qx3IVykucaHXTr2l/tw610d4dEqneAPDGA0iUjvLSRWGXcpVPtD5LTrOLXPhe01r+Wo+qCq6NVtElpLMn78+DER0cDdcaI8MZ/ORGzUSaQrtGLzt69r08Tg5HL0pLD3hXyu3OpV+EvHZlCtUNDM/5yFl1mggiyzwEwSXRHDxHc2QTPrnKe0mZkHx4EoUFuzyCoQ+MCjQO1TOCg4Gbzg7R9BaUqevEx0irX7v1C5W0QS4GM11lZejk4RJYe0BPkAAGzpe4j1q2v3mTCvA71GWW3vAHrdEDvBwNVi70QtjJQ4UXwy+JVedWKluli3WO75Nrrihj3RnowDKwiceJKTRKhp0rEoYx2jZ5liGgd/gjPXkYOGWD2lO5FbuQDlNcveCQSFUbGBs5YyG69auwxR8JEKCg7OXF71BN5YaTNKvcEAEbezgzrOvLFz8oKUxkLyYV4hMPDEKpNRY8dZlAMUrlVnP2o2iyuFsDIdEYvSJWvGsB5qHEqwgezLHWVdXUf8x1jy2pQDZqqvlivlTgAxSlHZMAcnKu8qo013Irhvi+iL8ASgvdoQ1osL6nmYZgFpdDL3h7NYSxicwi1NAS7zX5YHOeHywt44F3Oi0vxC2MaFzotC9XiPPJGKbQrzwwDFrVWybnrtLKBhQmujJ3qLCrGXPU48FhLBwqUvMZeW08bsMm8Ou2V6X+INFYaVfUtjTADbHUKjw8zVbyTaauNVmYxgDtTeopoLquIU6TIHVfAkalnqx/k8XBqxuLpQXU1/ikxKeoADvGdgfyL+Bju0ncERNjQ8HSXQ7GtSZyrnkjzw3ozaqKZDXzLMI8Hlc+5lz+xH7pIS7/RT9ylyhJDj/cPDn6HgFrF9Itq2ci48jtKHCXaeilKTi462KaKYu/D4lVguDVCvTRqIYrGt/fdDxcRCTRmOE1PMALQ4OPwECgCB6MowmMgPUY8ki22fE51fwD3icokK2Up39o4szqUiaOeGW+2ZpHOrkw4fEwk2t/fQPcPMS7QGBTETJrpW+Ds58sOgliAO8V2Cq5V56+DL591vo4/iQ2ILW0Jk13M+8Djn5FDYlhxUp/LfarIHyRefGcm6aHgRviioXa4NUmvXMGFqZneXUZmTMFhXBqXtDVnKx3DLzUrdQDNehjy2yg2vZXm59mHixoCuGkto08wHqVS6QWfB7zNBgqABgeScX4l3Gcl+hPtQsVZYjhJ0JND9w081K4eOwp2/pB60ra+r9KhdUKI+1Gj13iOKQl1o4aeUrMC2QLDHDyHCCcwUwbu1rTqe/e9Tl9Gxy3RDINalBEDPhtJ1MPed9KpOix4Jqgcah1Od+0OXSFqcY6e3aMazDEra3lnepgUeHLyJpHK8RayMz1hFoclkpTTOpONQjU/3EvtzLlIwWdwJ8B3iW0DbiOiM+TA5NQfatfmXKiS3YpGYOpFyS05t5w+1woEFnGtc+Oq99JZnVakd0F7kP5thB8wU/WjO5gHgFHIuPLxM2KrR9DD2haQGK/Lik7kxf5Uql0tV07NStCVF0XVZPDNLTtZdAg3NWy0Xgf7F1BkQD3h84hzD6Fs9uAMdXjwHvCjZrLPkh/U49F6hhmD4RD26cnll4fajXyXXZ8RyPNKFHI19yPD1vUvFOviGzAtxhNBLLY35PBjV6iXVcfxJygjGvd1Z/xI6qgRE48YJzBBEpW3lt08QnNdoegp2SyXsZvUX1LICJ9UM6r4E7QLnJYhHI38Qem276HFdPKSsZntDkB7AwWWUFYcImPuIR0uBe/A5supiLSD8kVgm8+uh8gwlDWhA6NXiu0sxpuFjkQ/NTLVYLvph+Vl9r8faJy8do1QLGfrGfaYY1H81JlxXfJG7KGdxgVHy1y+pZLe7ouRxrT6JWE1DIXjSeyy9HlyO4vT0IxXCsO+t2vVzH/kLCeQuO7CJ4qi+tqMyorrMSJlFj4jmC20E6tv2j4s7UNyuw7jUD2jzQL/AIO5Ncz3VDSsD3cMN4gpHwKI0Asgd2ac3rpAFHlFvlMrNMQUNUhY+I5cNuQdW14CJiBbNtcpd7XK2PcCjNd1briAsufHMacWgLlj8JOPUBKZbEA/9EeCU9zk7hPLAjSyY4RJEfDFAt3R87AeRBkieQdTQrXzLeraYt2YvQoVnMFcAr2Rlby+WWuhZUvlxo7dO8v72tvdWNiBLKVOdxdVlKdAjbNycfMPrjobwrHZrpEMAbAq0Wua+IVDgCgGl1jue0JlWBDwS8o+HIu2jpp3uGmlQzCNAYQQPeHKfbTxAYZnuhYnUdTxEQ7TwBdCw92K7gOgwA4zh10g8rAvDofghOADQDEBIZG1rwMEWEy7O7u2XtKnA3Glmh4DcgMhKDd9O1NJ7we3xGCVTfvcOLpgBWYMGmhNxEe9zcsQGNI+NALq9dqmWTBt2atxBCOuDoH8gEmHg1T2kvmLgsYNKwaKdzaDJOLrewDdmiQgomiVFZqhU2WeBhPMCiuz9aTRMXXvGrqfiVrYcTNZ5Kx5DGO4YzaQGTT5lHPD+JYjh7QOEBQGCDXWBaXTd2jsx+h2W1jjg4fMewy2tbQZfbgO/LgP5Ixv5q3qrOzF1AQZrCEq7bBHWoPVc3xc2v4xDCWGhHqs3g/sZ3muwOWwf7EUh3Sqdabai9M0yhs8JY9GJE7NZ3JiNeEWFImsHFjNit95RYZsl9S794egiKMeYwa1qB2YsSqYv+3VtKMOUIfDh6xCvAOXgR3+kCxhUmrINbXBdRyZwu6Vla2W2QRkMUw6ViBWld4GswEhKQsTrANBBB97I2+IGsUqt71s7nzAmHobPIZO4+0oFrVNooyihfWHWnVIfR1e2I+CSxyGCtfmAVpcr4NYcorc5dr5JQAjVvxXVPDTP9poD07WOsbiW4YXUVbWjvCNlFb9x7wMRCzUJ3gGr5lHQuCLNekb1eSwOuM+YmrCF+JZxxcTa4FzXuH69pV4+DjxcFd4DSCmd6Up8wsgsZT3gWtXEu194AcU8EOqZAA7aiGgja1X2feJKGwbHkEVYUs0ybC0va4IYtiHozNBIYV5lFbflnQ9kHKynuyxAOrCKqWjqQ+ZrVgEt9xlq4joh7RUajFKPtneqYIUZ00+IniFpACWFyssPujzzAaKTgR29Q94QErUoCKF4RXrDuqAgDmmsxglMMVTUiYhszc7Z+pprgS34eEy7SwIrDvkiuntBCIGW2EUMFBtdCWNnh5bFbRCenlLXFg2Jk6wiHyqV+5X8OTL9Y+WUGHaNNB7S91/UBlAZXQeY6NqjvaX1T2mqA0Vy/BbpbCIDr0qcSuCgLRwVuy4i1feE8DpCrxSUHAQHHtpL3WUjenbEvTffDfbf8JeTN92A6rkXpDViudWtiLtQnvC7zFrvEChxrldia9ZK53SbsIyrEsJXOrNkD05bcSqNTS6QzqALzcEYgViCfOBX2cxUoAC1PmEXjVcnUPbeUxrLDHvSolS06VWhfLp7yu9ohm0s8CLchOqXDqGPbXxLzD1yqtwBw14W/A1l8egJSZEqVVAdmf0PMPePWa4onJBFXW0s5Qv1inQ7rHBktQb5rs1GFiKOALDOmNYOyDiL7SXsKvxKYcGeS6/UMOJWImiiWB2/wBiK0xq0XFaH23geCF3Nw6NoSEja46C3gNX5lirRh5KfllRMYguCwHRIebUktLsqtcR9HQZ0vJ7TAtAFkM15gWS/qKhkBtALxw6lunh/JDvBmbkQzxgEuhzWnaVK0uXD7wtOU3I/p+O0JLLgKLUeGI8L+cIQ+57R9xMLdarl46TSmyaCVL9gtbAPJLI4tqm0dcdoqkgxwX3/wCRXElqgYtHqBLCNhxF2RNRVjpLxJ3uBsXutnaAmBY6GHhHzhgIUUjoxTRVicbnLjtHRdopQ4S8kHWQcK9HJ+N5cy+sQDzGjRtAJHZRGx/ntLC8ix56yrpUMFMHJiYuGgK8m50YBssgB75sZlWIKhWyGcNNntAjaKJY01s1OsHYQclWlO3NS6XF6XQSdv8AMVtrAqqHWajAdRhwqnBu6n+I8dfA2a2X7GaZPkA7Nn+pudr2adSpgiyyC3VoIUps85ZoDT2iU28QA4qM2xgQPLivKEzPbvJWl8XCBXUFU9ab9mXT0yyHZJ/IDLKFRYYe7CldZIHiAoNs2CTKjM18ZH+aV1hd1Xoq8DMQTEU7BfKWsGMqXdKrvFbX1Srmfev1GBVB1N8F7l2WvEtIRVjY71qPTStZYlVtRdGU7xjjkiPWskaGxQk3rA9sMqGMNa9V1fM06h3DDWhXJOYL0wxBR8uieZRqZyrru7FsRrjI1gtvHGYHmgH6i1Yg/wCiE8rUip61AQ5RVp3v3RIVBsxR/wCDMaWhxD5Hwy2RZfLP15jFqrQznLZjq0R8ZA12MslGMxEo3sOxFHeB1A2h3Ttn4hMyznm6Oh6iwMmO2k0BrzFrLnriE55VVvQG7HWDI4ewy9jzGguhQI5Bajw8sKG+RANHc6ta4mixKKumGXpAo+007/4jFnTBFPC5Iga36yzW6hsDWpoCLVG3dS+neFfEC0tqJg8rl4iUD65A2Z7iqu/EzAWiAJ1LQ9odjYdNejrACQeRf5HsgF1wuRcJqPRio+kDt3gigNA9m+OZR+VyIpbzu+IDlJKkWNSjAWsmWJ40A9BCMKvG0coSi6vtCrEKy6mgWb44hbH4HJ11PmdYL8LKQ6Rc7yxTzN12A3ViasiVGlodsHdJjF1Z0gOWNEiA3Pt+mW1ymO3bHq8rZLGXKUC3Y7wH3TOvDpzVlOsvhy2s9N7pSHXosSxJePzFc9URbK8fqHcCA2olly2WP2DsW9JYHmqtlD2F+EYNkBMm2iv5lLowmjdb3MGkEEWmVuQ6tdzHSLQWBjv6PjnpBFmZUKyg+jeGRhe44RabRBFaXrhHL/TZgEyciwWUMW0CBcpZnNuC77vd4RmEcddShu3b1nb/ACBxu9vdG/yPdFt1LIFbbQ71Z8y9NculfsI1zP1+rgtDq0SgcreiuB07e6BjkGsDApymB8xmd+lYB7GIoha6IoFpl00zmGBt9Q+ljvy6Qk8YV5W4mo9GKPuK4EUfGviFtPNoiWMCAVq0BDC0cryKdX0MdYxQ1DA6miPnrBYqt0W6bamj2i/cw8VzglyYWXCO7jJzfxL04HEJSdUO6zrGBAykK3SE3E8kBiULi+D0fzFhxLenhG34DK9CWU/avptAetsFkmXxTebIUDf2Vvy5IrjKWiaFbNfeJHcuV2ytpy0McOdlH2aR5U9JgwMkInHBfxBhMIWE6QQMtHtLh1oa+q0HVjfS2xYjjU7CiXFowCP2ckRNDCDyJ8JjWFRRC7UVdD3hKvyzc+NHUjasCkG8vM7kzxUUCdtzrBepyQQkWpgJWdnJdju9PdByewKX2ju5lb53Q7BNe+sNRRlsaoYZXrCxrplqh2eSAMpS85XuuxghSANHoTELZtqoneaV/MLiwyW+Ayss+kXgC09DMLqtQau6u71YGelbVHahL/Mf7AtCVYrjpCDtUWWzydNOkvVKbQ70/wCoPpIMYONUdCpkFCbSRX3Wg6s3z0JEcavYUQCJKqQeI2WNijewV4lfQCJnWqe9QsICxDmtH89ZWGuFL8zU+ZlNMinvGpbvygQDWq0BLTwy7XXe9C4Y6lOz8vdmX8yFNKmaQ2uToLh6k/4H+x0iK1UK3ZptUa3ajU8BaJH0KO60Ch8yuc6Bb7RMBA4zQYfeXgE2ejj4nJDYkqgn4j1IqPUuoks9dgfBYw9KGf3vOKY7V08UrD1SWU+iGbGl7EB7wi8lazkPM1C8EfPR6y0Atd0j59zvLkMYt/zhOpiEDBaiPbmJh0inDlUr8orBCQ2VyyDBTwyhxV/iUUgD7nOtdtYIuKDD/YKF46zeX2UOQyPZnVhSHTOgOtPeN1osOvFkYfe8bFas07Q15oI3KWv05hFkFrPuUMHQB3leOUVmXFpBjtyCFOmsGplUQEDiYn6NG8Gp0bI7pmMD5PXv7JYoBpB2cwgjbDZqxqrpHwamW6P7h5YO3qmm2+TV5VxVQLUWvzNUprNyW+7eDwGAoBpLK1c1Cwurt03uTW/gRb537kxpik8hNg3lox8L+2eA2FvSCoZVWTjeOp4lZwVxykGSsqvtDGKBwJpdfMI2A7DCxbAoaBoQRqIKyXHWvTWPYO9GWuhoD1gcnZII/TIs5ej5jEYlVDJ6qLgKDDUbxyv3FeA6BRpCwmCLHYUvJftGOnt/qBgpHcQ7eHOfDMhzCrTRgnCQc19regeq7WdJfWjQYaCxbEIJa8EnOMBrloh+YIx2lOdODuwzMUEEEhy0GTr0qGKhsReyr7GYfJgXwluS0mwltlYnO7JU8nD1JddBQur8PdLNNokgMb75GBxGY7hdBZwPM0sQKf2Du29YlYjEBqwbdyfxEMMOwCr3DXugaiXNs7zVd6JFdzKg3kcn4gC8WgJ4++j0iKl/FldOqwhutdA9mO5t6TnZnreVyyrBpFQEIp0OuA3moDVYy/HNBRm4nmCisXnaAUDHI6nvMW7QQizQHvnqQNqp1RpqHuY1l/8A7SFq0VaQgNlu/l13x0hXNAdAdCVZ4jlhBKJrZdz5CAkJivw1lN8NhQ7q3RIXCUGrysDyKVyS0qm7J1vfefYy1TqES0FhW1gkqVy3uFuBlHgg0YbE6aR6EFoK6wm8Slw4F4WHHyRyNYCbJNQyl8QP4dxKA2X0vs6nDLk4MV+rmu8dSabEmRN1uTziOtnEOxzpL0z1mQCb135TK94RoDqykpDh5WiuyJkYtUxtS6bDF6lad9ncdI6uuutwG+/5EsXtpnN6FDO6YeIwRw0t56e8ymCxe96vvjpDZ3QqA7QBsEuL2msxANOpwxhtiphdcKdSCAaG1r1lXqwpIGmGnvmBbzgA41uTAYVuQyYW/HWMgdkWdNg6EMOLmBVHaXYoIWLqIBwjAwKWY/RdPOI3zHJRyz8Iu1wsGHkxGvbVsTY6/EWGymCzi2/37RE8WqPlMr3hhQ+CNNyZrCusDyVIkThIbAEK7cWWuozCX0S1yHPZBlWWUFcdxo+TzClOZEB5v/YcZWzwFmezSHl2qQDtFigWE1VeJrtydH4iIdETQhpnCYIbowspRtghBg3zBBTHMXQOhgJhe+GxQTWyaaWqy/L+rMuym1Zri27a43xWfI5xQQ5GEBLHbQx6rKD/AEBfV1GVryOSDgrolKGnhgOz1EESC1Kohp7aVOwMr2xE6Uzgq7DEihPjUd+XqwYalHZsxl2iQMll7jR2luUuBu8M1CLW9OppBOIigOrDhKIKHgrU6setNVX72VdJuMgqG14exFnJQ1OrsOsOVShXbFy9Y7lggNCMPHWWf0iF/K68dWKNH0mt7eLmcCVAu1jpGCbxher/AFDv2/7LApGesc4/KD3MAoBoEq1u7wbrrqSxv5gJwK+zBEpiorpR4DMUciAhUxDKO8/UvN5UdV3uXIWWw3lgUTkBbuurKxS3dgrga1rAbXHbWGUInj3RwRXdUNpTTXYYVAoKKjKHhq7X3Unll1yktXuy8Y1mX4qNfgLTIJ8R+ZSDGq/ssuW6TmWWEe6/EZjBsJpo8QEqYDYCiENXBlhlOxTJRtwED9DQld800xzE4jLQmC0K1d5YSqpB1EASb2q6l+zMPkuG5CsDEEJOG2emLKxilKxXkgeLmTjBox6UM53PuGWDmEUQThi2xhhSiwrOtxOtiTkSCyCY4y23FKGD8ivWDwyxlVjZCXrrUhLbkL4a94dY12lpcK0AcxvGXbq23hBlQIiXjNwFVUcGXMawc9a7emHOvvFpwK6v7E2zAoAVnayBaNYbkoRYmWmA/CwtDXKug8cwHwKKuyHPeA5nT948BVbi919H4jeCVFE8xMy7DdLOk1rODsn+7yjkVqhul97Q+I9K34fqoAnhFWJzcddIFGPLAN6yochrGOgJbB6OWnWXzQIBDzYxwQsDm24vX3lqlolkwpTUnBKiGMV/cAwwpWJ3l07HeZbeWCJUxDlBais6NnqTXGcBTytEhhOw1w7irzrLphSXuZpfdMC8GR6ZNn4glCsWxO8UOEXG8CmlvKy67z0mLrEBcxqdQ6j2ly9qoBdHT8pYUxC3Q0yhVGO6BJEFsLUeU3Qz82ID3i9YDrBBi2WaodJlUx1hw8yITtL1S6Nt12eJTxLPYYB8o9QVNYjqlj5hWNMlnz/EAqReekUtE0VKRzOt94gmU1QoKV1IBkDD2gGtqCIlpYmsbmOjIO7tLPOJQV9No6bDJ3jA2x/jIdEVTR3h8mRk11X+JvCyCSi5Qdb8MPUU8kQXsFIZ6sbLHDbXrx5hl+DgE6VaYqXpWe8KjoNy62Qkm8reO6xGvURO6dXTSHZ+h0BwEGtlMDcmOSdvkljQJxGQtFYgLqFnkI2w901BVHKOXscTjx3ZgNoNJ4Jkuhz0Q9bE1C9XY6ExLLIIc9IWHwyvd/CFmEb9twN5XiwES2wui+viL+Fxtq1doUQ41AFc4PzK1V4H/ZbVpvk3Z/1DHxACgNggjBUx5K6kdtZyRYjkVLwHK8Sya+Le6V5d5ZB6QN7ByioctYjg6N4f4OZ8NyjBnSXIYWDG5wBuyogx9G5AmoRTudoZL7ppPzFMnxwDK3LTRmGlwd1ywSsyhRQq+JfXYWCLsN9JbzNNJTen38wUH4UqtTcRpQwmi3mWEOForZVbSg47RV0dI7XY8k6jkoG1vvbzKBK+RvDAAWq4CM1dBFDoKIGotwKywPxCWDS3dENTLV63GQh22lEQa0HiEwiJhmpC3ArLt8uSeePE350xvQb7wMMOCCOA3VYtFSqAAZWwl1tKLtVpVcqL3WZXqcfyaYOETVNnTTGGVTE6ExAgKM2rPzBcCCL5GudVA4lwjFggElq7AyvaADnI9F5dC86S3m9lae+qDehvqg9VvjXxHaQsdeCHfGvSat0D4j51Ehmv2k2Dx0lhycn4hxx2nD8Q6YkcZdQ9tAPll/AbhY63LWAPSR/KOkItedO/eWzLOnXA7UHLPeWXr7Wx9EWHAi1PW7ufiCzGe0KrTMFNIAWwBqxEEKKh0YX4Om8WHlhaPMJAJReN0OfZlfoL2NGVd23xK5zYy4iaw3HMdoDCF+F+iPpEIq7OZRqeWAJpcCn6iKlyBW2672mfWEgJdu5/A5jClpBH3lB3XIo989HtKpYjtVp6Q5QLw4lfO2ge4MnSc3mQHhNnpLa0pyyxKvwQ0lw2YmUBFqHqWzGx7w2dYMFaLr0hyWQf3JkJ+BUcbCniPN6Gaxw4bHJC5cI6OpydSUGq+Jhk+0eJ5YC0tgjdDHWko1tgVl0jGoW+pmrRdImhbEntYVKwolvnak095THTj0MaGy285CoEXIRr+x1JxncxECVaSzQSorFFI2PeCMRbtd4h3xGG1VFHFFX2xFFbLFruWLfmZEHsUgFt6NtpSeqrP3G86Kbw+hzFxuHfEQB1IZVla1D10EJ5hBVZtu9oIMaJAUxa0Z6aQhU2pZzdveOk3HfcL12YmsWoK3U56xL4MeK1zWzqYhDIDXECYA6M2HqTiD0lQ83YL5dA7xXadSW8hu9XxGzyPnQtcVTUpSkpFMaABCstusOq/wCIMLnEXuMaMxCNM/3H4pQGrOSUBVdEEVPcg4CZQ4JsKbG/rscQLTg1wcPxGe0GrORNjTDXqtzHAIFLyux3iCg6E2hZerG3f+Kr2GYdAdn3PyE3BCnFWck2qLw4mh6wbPLx1RaZoV78KS3l94GNmYZwfOxxG4ZCJLYNVguq0gqdKyr5gzBcLYNFuvLDdzK0m7+WYd4ccJFb7bnCYgARy9oFqV1hBGKgA3ZTODTHNPxxCQPlDBn81oR9BGNCRtzlz7VFFFGqjquvWJwaZCrtrGQuKlKY/qGGOVx91/Fo9JdpTs6P2aMJY25mvcd9ImiiVAJ+Vy9IGAWGFrWNHZbMVzzLDjMuzlkHoB0uoBwxoICOdZan5FN0DH6s8/YOHLXUgWKuCdS2rqx2j591FyisjLPHEERohulwfJI7EtYxXOfEU+EVlcqDdzoQYwzIDtc0XHzGniBTrAZVtfmA9Os5f9IXitMOHTfKynWpriVYsZ2mJjyihy3S554YnMYawm6MicMRTx7zOik0cUNHbLLm5OvaOIem6IMv4gymYpwLP1HWKkQpXmgAniaBxVhWZKPOOPDj4kIQ2SAEb+YnSbNr6ZuPGjrCMtar8dHoxNLDPIhCdKerhYa6auJfZESts4i+E6asCksmML4Trq7zAcqTJsGthw3DA9yXamqIovtwv4WK+qQ4RLpJXXPc6gJpNjPMISsKZEtCMKvstQrnWmHHmUT8sJulqUBHjObwPIur2HWN2D3/ACSsrKnhoyhwtez4iMFNRJgjTXelYVHDwgug7OzUp8aiKXB2OGeY7ZDMq6hrZ3iCAgKivU6OpFf8QTStIAmaUsdH6bvzqwz+USgg0FphwmmNm3MTOqlXDMRi00DzGrv1SZ+oK/5HCQKChWKdTj3xTywBvSLm3ztESB2Nse0d6/xBjPGVtA1V4lZal1AbKNDo8wgEh6BxUAlSXoD3SOjmqGDlXkiJmkKpm8Z5mfQwVcgx+UJviidDHyVKqSa1Vbl6nWFHKEabrHMIIxeUO2x1cQr91HaU+ZhOkFAELqCGXh7nRg5bLvfplh7y8obAO1oX5io+odO+L1dNI6EQTp+l+SEXCwFiM+kjEsU4j6iat/UHzBKMoWD2HfWGgFdpiSjE+F2jyKtgjhQvxChd0CPUP0iu/QB9pVeIdnFGAP75zCe5jUOibRi4T1YnSBrULsPySt3oQH83l9h8BABo6Q+ysDo9LjUi1ZlbNCXLSxU4fAiiPWf8RCsl1dG2F2hUZGRhXV1ZYahaZF2ISSTa1pbF9rqD7MvGDa1tVEozYK71qLeRqBoUmaNT3u+50cQhVRNcZ/zQAJ8i2MMBtnl6BvEkzrv/AMPzCSSKs8lXQ6sTOPsWBWrmU7tKQHQGCG7ABO6u7EaGIkYLj2hXPCIfiInZKBxh+bRlaJLGsjJgbDK0BuyppAHU3RdnEr4RaA9VS2VF7th77YOlw6MqGt9DL0hlPyuz32OkR79ZUhTP2HUB/TiU2GDXEf8AGwsZNKyPF1g7u6/UF5WFI2ox3IkGokbGD+Y3W/XHfsQRa5uL2mHZKXuD5YLtEUaTIABNjjo6OIsS6yuO/wAT4hYACiKCB/66IHVrZtzCeYmQXV1XjVj+pBxDhR7wEADYircmkYbFbDljsbTJ2xIbKhL6/QGnQZZ/lP3k1dUr1BBoug8wQYSRvTCZa2CCDXlXdO9wZgI4SYK5xMbhY1ox4CoCZ2M9yYQb9vMJiAbQBQQqauAJmw8HjfMbSiCMXY/ppyTQHNwVwZ93iM7spaUoXYOYGJsKiUrk6swpgZdXKNjjCrDDXxEu6MpA5eIfWVrG8F1q0hGeOGMiY8KxEZIHvgFl7rsyTBY8/hbHzzMvilRbENN9NZZ4YN4wR36MwOM0HI8DpHmBgi3+vDuH0SOiG/MWpxo4lFAavchmW2gEHQ9JhWJHqDbmtg2DB5mG3LC2OBBpOIB0yQUxlzApy6g5Ade7HECis7g2oWaZrCAuh8ONVlomjtEXUQbxkHRpekb4DotviXBlNBbJrikJxWeKHbdLCJBS87z+UYmAiZVk4HU4SWjZJoTA1cHzLqTpNDso0OjzBTKB0BwegE5PRkSJ88OCOov2e0XpFEiCmR04xIARrTMfZ694BAy55P8AhNGVkTXl3LNNiCwy46mCjRlbdtF8b/zEIBgxRtC0m00uVZq6Lo2vyQOh3gCiBxTKHAlOTDjdbks3eOtu7NeiGSbjK9A5/SK0ENB9gDmKZOdj+i3MKjBUBhumdprlCwvuanSKL22jyj+Rc6nKIxpg+HIJnvBR5JU6LX2agFcdRVzfsTQwQuPl5eCZ2/5/SPwEY1gqDWjTMJUGMaDYkNCOQmu+/iVkhDWOTmW5RUKeoNgp1giTcC+y3dSULEgPJwuYE0MxPbNwbvXQl6KtryzqLKGQI0cRaeWIbaadYSiqkNm11r5lnkGngWlr8QY7hS8IhTNTsLonZg/dwKnQr+S0/Xngdjr7QCOsrVd1d2WTVHEtqLF73rDtjrN70KDPqP8AZhHIc1p9o/lBFqatqVwYAekAfIsz4gtw9UX5iZDmchmVtLOJTO7iBkOpEDUCTCXKEbA+R17tNmWAdusuguh2hq3UFNdUMsuH9QtnKQ8JnT1Z7CrX5jXpRFq3SG0eJWuGAFHyRQWAxEikIN3AWrhpoXZMBM1ao6CLkN4yAVdrDhrBrIRbqKqqy/PNGAdbbE0ri2HggcZ1mW0qIG4lL0nE7Ry3g1iQd1ZSnh6HU5hXzh75eXEKl2BCucCwEUkhQGE94F2aFd3p1lJH29R0j53gLbKzTEoZaTGpoa8kQmqvYnMY6FaV5WbK11lgDUhVGRrWmB0UzE2rzvweZRVy2115gcIKY3RmxsaNX8QEyBqAbE4Ewf2Gj+GXjo2dM3e1cxwG3JBVvjeM9rjl02BTN6wOFRLuAoaq2/f2ik+t7TNWgLsxfEYG0npJr5W+CXw0sYEYlMa1RrDXNHUTmZgAjo0ZbNPzHuR94+UgcWDYTcgAGkqP+URoCq13vaD1MAjRVow9pSJWamwbTDEKNX4BBj0CoNcGsXVDTNPiMfbCy6SzVcF8R7yAV3bJT0OJ8lfzRDj+1xwOKQmI5OR7qaQShpOYSa9YtBhWbMOgvVe8EsnFoC6s2lGTg4w2NalbdYU4aBQHQmOipgqV0ZBK9FqR0b8RGschb0RVzEayOAH5lWwRFbH3iwNXOmL36+YnORyA3GUrNupDqHXlmmNrdL6wKYroSqVpNeUsCg2jZ+Q5O0IXYPq5qh+0ZNHhQ2q6JMjdKdUarqMRAA5hcrruEIFr3KcBwRRBQjE3gqB/sNIoi5Si7JpmF1tv3fEqant/U2D5B+pqbEHF9ROXxL92VhrNHNn6EPF6qLoH0xKDhEW7OSNzToyy+0rOJQq6gbRoaB2nHBnyiC3wdmAmNpx2TD8MeB4j9SnuZjT7xLRrb9YU0iklkEAKqvuOsMiykA9YuDugpnXpKCwx1llj8Slf3F4oF5h4CYSr0m/IaXWHowRQO2JghwOcjUzaaX4KDtbfNN8uWoeE1GAhRHMy1agZA94XhzDDvcvQJqJYw3K861G+h3JenQIvJto/EcmFNcHNpme7a2a68+ZaZ3Yx5NT5IGUi7LGLGBFW1xeiV4oevpAfxKAOZ5cvtCldUby1mVNcza5l7dBAHDHMdFoOI7K2mHjZwh6sSTb2B0P7DSmgNsb5JcrYgOucGXlZZBOGD4vwQR4YEB2mLMIl5nB7RGi7Sigs5IcHrpgiQYhVTubB5l840i9qWWhAuQn2Kw0e8codOl/neC9QCz/2OdI+ztBopmXF+6dCcQ73uUFksnQDVWXJXg9/hOsBVfidjlFq66xAIJKO93tweJrzDikNGqgKjdehCxw7SnNmh+ZmMY0gVOhOzAtn8Uro04bxLFtwHKfl8SqHTwcDzHwiTujVoc8p1i5LMsrAMghW6m7A1XQIR8tDVdVMV1McwMFkZGsNa3gkYd87MHf8JmK6A0s+Z1hlTMLXPHxAjmlbuhEd1ryrNAjA9GrUctvofMB0QugFEApBXSaSASkFeep8o72qIoUAexEVFo7mkK3tf4YAmDJtdulnY+YgNzZswIhhS3seucYgVbhYSxaejQ5lj00mKklRHStooZMtoDgvtgq2fltHnG0jeyJriYZRBUcg4Bu76wbCHSFZJEzOAKD0rnvB9jEeC1mtNYTU02mnXSvzNeGCOzfgt8RNJo8XdfNQq79CWrenEFlQ5Mw8lQ+mnQ0NC0s3ioPSFnsXrpEkXyht9o9GIncpg6onaYTalb7tEfk+24b9jZ4m8NVowe7XzNAnzLRQl5nSZU1HCMIG0mA10v3mskymr8WHTAinYduzKl9gXbh0aBfMvTZZ1Tltw7Q7QmhKWB7mjA/Ihk5JkyTAxu5DrA6kZAF3Czm+GXQC9yW+fkSzhZdX2vUt7TPlssi2O+u8zGheFXVP1UFxe7bE5ihEDHJECmzeL1ekww0jTtcOtMxpoCrEYmHZCd7nqijCDUoSI6FkK90ODH2z9kR8wiMCZVbjga2gvUdjok2iNlDlMOrfT0jRRlYV1mdNZwIVCtUeTudNYtgtXeBtQzAvNSomlU/cGWM1ymo6PeCWnUP3HRiLzBlTiDWxS29NZU0F94GTrxBW9iaIuGGqrIYM60aN72OzBHyAtXORPM10ECD1EjhHI1HubzbRGVt77eY7OhhG7hjrYJYc1FAwV6L8UgMtGbCQ1jSY9bcxW5DIy4LOb2MwLPSOtksE28xoNzSrL3/iA2gIR75YlrmCLwbvzEaGJ382K71QMQiw810OhLDBnaE2plGEanBmZxgbMoTSQCf0csCAHZKt03OjvKjWZMA621HXeABkoWjShweYs4OwYI0qRfc7iG+lTFKbtuggiPYVXWGqO4mRY6IWr6DAtDttiVlIWxfWrrvR2YUQWPJXqA7OYVqlnrxVtYga8chdRoJ7ux1j1AExzju7JLWVoOGU146zWiytSP8ABbyor5m1sdXxHwiVQQEsOmrliAt0WmY5Roa0uLjKlY2Be05y9ERXdAbsm+NTELh9Ij71AQgFgzcCuJS12RV06yy+3GpaDqsetzAFjj6GPabhY229BPgJlwGKJdb4WFOIzrog5StuGh5hl2PCLDVlpo7u0zInGkbRz4NsS1TXPTa7Z/MEaigsw8QlDg50ZjXyzbzN+B7wARDYGRRiZ61WoGwX1Pcl+uUa0nqLgBHBdNoNMU9cfMVlHBe+Yw3KZUeOAQ3hJZC8qWsgEQhG1O6VbQ7+ROpOJWrbrKbvuAclH2PMwRmDsU7DdUb1FY3E7vmp7Rli0RXoKt8u0rfiEZYv6R3QKgatj2w1LmHKgHvGpfB0g0FhPT2cyjmrdkKUO4V6jrBlLaWKhtK5ICxH5qAwEswvUBxkhtVUmuBbyX5iFVN1warE2VfLxuZY66yAzZssdICvDYmG9GneCjnaRNtE3q3D3Ljx9YV3L7LmawIgHc3v8ygA2a6/5NMbxNVc7VDw/BDY+TAtwXAd4AfWrB34T86R+FDmk0WxV0Nqhye1Z7QZ/I4AbvfFUoaAAF3kW+CUo3gAI5KMD8x8xUED21EwyxdBYneXTjpAotwiXmd24UqAyroQlgJBCbyYXGdkq+kpEp0NkCfkuNN5uly7Zk2l3ubLsdSoGGyNz3qDb1uFqpGiL1P+JW0lhbRFC8jaAjo6LKlBDad0veEB6SowtWHW9lGhCIBw6vVeD10jaDBgYC5N8KYEqpCsyOaX0hELWEA0R33gRQhxW44vXRlIDlRbm3SUIwJUyrjtKIo0tr0A/e0RLhSAjamvKLUiiqOh+YSNmxd+VEtk4uv4YY94aCKhO57hwzOO7IN1z747wJTV4Xg3OpGzgt5llXiOWJR3iX6IViJkddBU46XEVeyh+yDwzMUZjE4LBgpvRgoO6yQgJLhJrjX2jMOGBGBt9jbfmVSaVX9HyJ/w0ybk/dhsYj2I5B1q32DeJ7zmfg4dj3itnoimd+XVp3R/IdorvJ1esZcTRa+a/ZA7hzMHJ2yr10IN3rg6EuFKnGJomyRQIe1G3F+cIqkSxgaaRoaXA0tLxCy4mVp05Y1sAUbLRcAOPiLakIWjTCoEwtrerWW1vpLmGUGu8AEWUqxjejvO0W03jErxWkEMwIX/ACfA2lm8B2ETYmOYllUgZiW0GJ5RcEXoiZb2PPV7RIIEve1sGDxBFDChAaFAQL6HxDo8KZ7qrBGIs0ITgrQI7kWxanHu7kzlsRwrtz4gKzk5iI9lBV5CLnLKz6LBKWQB7NybihljY2KxW3gDKQ7lWxKKzfTiC2u8KghoStcpuG8Rxu2I2qZV1EsOF34OpBJCL2I6JFRpOhgFoDpC9VcgrC9TR7wraq+ugaPYEs9XbkOxbqwOLgZ9tKG0FuKnQvH+xOPfP9lT5G0nUekQUsHUU/BnzARPrHPwb8aiaVKj8dNzhMMsa15GaBFx0BbmDT/wVrAdiiJrMEoK1iNb9asw+cCeUY5iMM3A9h94hQDgx/MW8IdLH5jMjKvCmKs25vSFkxPHRsa3NLlrUuhshzCIMslPbjeNNRE/kI7bS5gUeQ8RQLCBpZR3GnSVKEG7m+4I8Qa+FoFd33Zedpj1C3R+JM3HREVStXEoZmlXnUWrFSgRxY1RghSwzSXlmuEiQUHlhlLuwJtLZL037yyT9V0n2IUeIeRgBgvybwMJkAYAHnL3jpw4lqNys6Z/Ubx1rTWjVPwbQ7jKGPQTRbfaCLLrPPVO20aNlzX8FRD+bGWvsdUES+8xGLY1TfIxdC2Y3J6Hc8zetufK4j0wVtg48Dc7+xEfL3P4garDe13mnHDtHmChGFhRTNKnxynD+nzG5bWNU/7OGI0OoOVgAFHoy6XqOz3ghAkG1tM2zih3hsxUsaNnX8IBAHThMJAbreCEfDaKA6y/mCrZqu3L2SoHRKCB7FnLdgXuQV/yexRimz2mm5Xuipyc5kficQF2lsOyAIx0cr6MTAmLL4TmO9VvBFVAVqyma4otu3V7G0XApry9U3biAVjtFoXwieltSaFlhYeR3I2CrJGCBBN9hG0mXj2aDVoBfMoroLvuHXs+Ii4lhhRMjpNgA5hZdtW4Yccu0PC2DPDvy7wzCzaNTBKbIHojZl7ZfEUhK0CdLESKDxWxZrRljmixXtYWPWaApqj4dmCOpVUMOzfue0NsNpsYjkSyU5TXoSu3f6UaB+CCCAoBpNA14igR6kPitekeFZXRZjn9BU8hInUmf2eMF/T0dYuNwqKtvjadL8QuLhuMmzrVkEOlq0EOYUoIs8G/eK3mgcn7xKmd5tnzAxzQaPzLcaBKn6ZZQ2qlx41fiGGSgQAmResrYMVUHiDV1WyOyRce1Umz7cHeEAELNycumn4lcoGA/J+pdQGrteh0i/GwPFMPHgRDRCqbfa0BmATg5QoICTTH2ID5lumCLTlHAw4RMMQpvI56ls7u6Ck2ynI7ibJuQHdjhiti4LrHLwS0S2SrOht+UwssHVd4BWMQsOOKUPacvsIYkQFC3TYIV1qAfHQ6R8GajKDSJunTf2R3HWKOBgLufnUS8Vd32lSTUML1dCANbRQKoUNBenSXLARlvAC6NaEUGdlBLc6ynqeH9mSeT/cYH92Y9VTK1o8zyrusZLdYN50OxN7IisbO1rruejaBIgpYHeOWQmCKfD+YtSimILynK7Qk6CTMzVutb2j0YFT0/DXuyzH2eZavu+Yarg3RXXvLB4FGV8uIEgpoBULHaBioG8F3XOpH4vf98cmyRh8hrO/4geY8WNzG78pKyKNpRofwICFYDGAgU1LNtN+ISD3lLw4KIaNjmN+mBm4wmtY3QrRhgye0MsDqKspb1Fab4JfCbBbTHFtHeUuCrxeYdTQ7Q4QjVsdepWfEP+Zilm6cF7Qhw/K7q7rzCouhplmDuViL6rdnd0heWDy5o6NYSxLNX1yZ6SoxfSo/EosJhSKFwaiWJFcpp6G57flBlYZvbJbjbklaweulVD3D4iUWiy/hAcbyyio7qb7KugNo1BpMaaVVqze4q4/R2ul3mrPxwG9Nda8S25e0N/TNmFv9x7izyS+ydpRtE6SoLRp2nUHU2thOLpBH8hT4YWKu3yNA6csOsRPOsOMN3eNEtxWdmJYoKjOv+yCsSt2WEC2J2Ae0qQisaUTePBiebXQNr6aMtZkS5KpXJgvfEFGEcsuXDtDE2oUBHdH95RscdW8NFoygCaevEV28ymXLAf4OSW/vKsDZHcZTN+D/ABEan09pc3CLFjeyUyGNMA1JxFzzcU24FZe0Q0lYTiuZx1R5dscvY2lRbcrdqm6zFrEF58S5svEuTJjg/IsqGGxB9ww9ICX1jT+oLTy4jGBqw8xFXoWZsAcy+pZacPT+ozJQtGT+nWIAp1z9I5ZRZeFy/b26u8EgmdHzGl3MjxFCgybPKhrTkmekmnfSVskSkJ2RItBZrS9BjF8uEavqQQB2AvvG3cgXbM3D3bzQZ5w4n+CEiDQNIMqvxKW1mUsHELM+JVKDCVcgyS90FUg6wZWa43MwtR/2kMTh6/gm/DrLwQaBj2ftl9RpVMspwV6Fa+IaTLcjxQHepVYVHiRq6kFcCmuTld4rZgzJBaOOsO5CUgRezBD2ThngPMsbqmzEYzFOmOnB8x3xgvxDXJi2VeI0mLVwZg20BGOrqBOljLLfg6wOVL9Yrsg11gEHWLwWMsoeWhceh8XRjHiAVjO2oEp5dItOuRl2ejpFzEDma1HFuZXMJdQtA8Sk/PNWSupkkTpnuxuOkA1ntTK3abKQQO2XQdEljThCJopx3HJqXE8Fa6XANAaeZWaXWIZK9rWvEVdS6FuOGHDN9dYZrU6yRztCyvvCoYaFxNK7H5luZTNzXpCGCpC7I+dVaNraj8DSFAAjlNwA5d5VlmzBsdTnLBiMVg+B++xGkfzpOrrB/u/MbQ+/zNtI2tHroQH46RlGx7v4mAiVZmWF1U6CayXU9+iEZlM73YHUIOVwBSyTsWLUPSAqjaUOgh0YUHykTUAq5GVC/LhM4NAzm1YrWXfD2rHSqZhRw5uYUZLe8BcLD2e0C+eUfI7MrM+ewMUd3OO0rCt9mbHXEB2XN6ruruygxiYUiXTGgJLTR5fd0hHXGVTo2xrKsoqzWXI8Sj7FS/EtCsCslfoZ5oNJrzBTmT59nZMqDnGo/j4irG1rhHAbENlUs+ZeXAEFJO4lMqd4JqcYaqbxZiLQ00rcu2AQF4oTmfaaLWyERsguA8WiPDcVwv0wF+7mYkaEuAjRoBgV77UDQHPWEPU7t+00fzLhq4YRLHUY3Q5QV7OkWIuLylPaSb0OL6kq3191gjkht9dxvCQNr6K9BrrqJFCqQtDk7M82bQX0gdAdpj0gaxmXlOYbbeEvqdH4j5s5gJ4nL9XaX797/ELNsbMY1MqOELUdLhBCdYLqiahxKjQLNm5s73Bq3cNKZaXWULuAl1Kc9q9zkdmH7PwvboYeu8GgU0TL8TQXVkZDC1deYccjcm1jokmq/WkeGntoeHnmKRQcRGguUOuhG7piIc1M96QKqlIlj3jnlbpp3aPTSBZFxsS+ESNsZfSti+tQyNLS7zTyw5b8R+70196fMTBN3fvBAYygXQywYlhhk1iCZKb3nYWB2kzROGsPn0IawVJ0CLPCqUsQxMUgUyUBrzmBDiuibzhekAXVQDoDSCTTEw6Zh6MpcZgp1jRrRC9fadBEA2wjV7cHWP2JqXwlhbNlF1hQNRG27vqRhAluhsBeOPdUFeJHTWCZWhUBLd5cqyCm3JM0qr3I6BXWBqFHEAxA2al4DdioIgUhugy9UwksA1jcdI0zRsiuajqn6ukdRmefAv6j/o8qJf1ErSVhh04jo/CV0UlchR91gPVUaOo1uxM5SC6pt0GXicHNCbXAEF2XORG+coWPLLfbrGUaKFexMuCyVytlF5RlIlHzBrV2vOx5fglJZGsGnV1xZA5Gi2QgPeIsYyp3jwdo3R/D+xpVnj/YgqKzSN2VUUSHF+Xg/EKPpiAFE0MRKUeIAey3ohsUaMAiqsVZdlZDtLE3GiUanP8AsLTOGMMeEBht+an9l/CGRK7Z+InEQoOKboKykxLQ1Mm+UMIS9wWYaLiirhg51zqwQBQ1NyOFRFFcAeSBBNysoJbsRpQKx0TeLJZW2bFg1n4jm4cXwt0hkcLUP2QmZyYDvZ0zN1JorChyjvUCvNS5k0aqC7vSLbVAyv4iC+4FcFBMyj4HRHcKjCrbG5kdEPSAvjMQWQh6D5iuQJcq+kwGjTT+oZF/Yf7HfrGbB4PYXw+8Z2gyTnfgQ65Z1AJim+leY/wW6hFwnaAbQCjO+zG8zvPokGAWmSMe+kKVmd7DkhoB++sPynaWAksYtl2Tb9B0fDNAfTtWtLijMQIXZaPK6JL5QckdV2hYbHEEdvM6kucRqmGJeXkG1Hy4gKFOSibMYsjicuxyrL4TG+w90CDCJRbhGvQgBRKqvKPyICwh6xHNjFyPaoIKlN3rGrnSZ1awP+IFg4SI4hn3/FvVtEiuP/imsNOYAPqxAxkA/Mv0UFaackpi0U193k6wAAJYGxIhZZ4lKx3qLXDGxmHlmS6jjaVh8cMXvudGOkBnQ6A1RMMoKncq4HmrVYdYOMOiMOpNlGxOjR/MD2JZ9t56MAXTbzMrkwRGbu6j1ZCqiXDg9G3TQ6dXVmI5Vk9AuMAXAq9L8EEZ9OAdoBlLjvKpZtmXfMoLfJCk2l6h16HWOato0B057wFQVvEBNQaDyaBBNVJEJ4zEHBXyrwdYfIgl+CN3rEeJYFvMGbQOmnaKN1ccUomkvBVIu6N3XXpwdYShiwRboXHgC0K6DZUyOlVfglw58o/iUm/jHXNa8EW+vv8AfJFZhzLehcubylgU6GIogXgBvcahUYRyenBDKR3LXXHGPOkN/ITEb4axOab5Vn6hNFp3woz4Lly3gNOx5v8AEDyQwABxAoZiKwzTox2Vk2Y+1sDVtDquI0MpOLpQHAEKAOfYTHhAV7OZo19KfdjYvW0tM0T0f9jOEOi/sRrml7R4L5/EsptTcahKVo8xXU8DGEGlXaA3ZWCxOk3ezPeY4mr+hl+Ik4NzevJ0gRv1AafiX+ZHGs7fiBaoffeUERqH9opepndbvLFkWdX1sH5g8xxbLIAd6AjVSWzRkcVGR4QcfuPiNwbqqtXlYRoEHNAFQ0ABm1dF+DtCYKWDRIQoG+iUU27wD4YW7NKDYIQYygGGAWbkZBxygwt6RQ2CB/MpOCHwp+oUwfRfiJ9bYrMdIJq/xl1/UTMn18WaNS99otrC1ZycjzFU7vYyhhiACuJjnjIZgx7FAfImOalQitXnCZjrY9BITnwpBYDRrYHkWDuw2thkF8dILoOIZq/+vEqWWNjOH2czHhASjra2dIssFBZ3BNmWKzEy16QDogjTajr+pfLtrR0moYeJStIJZKtGMuIc20Vf02jLJB0Kl33MS2IEOJQ6HUvMFI5+wdEheXA4hTgLjW13gcRtJnpDJWZSht6m/MRUM8EzVDywQGN6QfGKJZ7ipmRek0apaxlrdcHqx05IH9F8B0SXSzCYSjLOTEyS14hIy2I6MEcqN0vn+PtDZQrKDEzNw0X8weaVgThRmZ0zZbJ0l3Yapw9Vs9NGDhOo3HqbTU0sq3EozdxOkizsQHaMaNIancgE4SW/LABT17dma9pSVwiRlbze9iaQSRcO5dSCFFuXhlzHRFvuNzoymZ4GicJtHQAZu9JZumrVk0dpnoLl+YIovK6FGmqr4zCbRoT7laRgBoZimhAjSpVNMRJyoNLL2L5hzloCgaodyIjZDVB4G710jYdtsL35jJC9XVznaJJ2Gc/Bc7deohtssgd5Ro46wBBAojbvQ6Qo0KJlLxKgiHa5Zq6eIrrAregS93edd1dpS85i5iuDqHRfq5dFZlVcW/iI6g4g6KjWdQp/sGRU7f7CpAjMDKCtYaEFTGTr+lXjaPsmUwwqCmSzmKtS+kBbWFqwSvxrj0kOETonGSOZ6mQaEB0u7YzRGgXo8EQ2g9BBG+5jPl1I03cxnqrgOrGwMwhdXu1HiHRMziZihcaSsHmMWU5QDVl/06BPpY4iH7oaUNDbPvUssdUYNQe7tM+JV4NdG7n2i2r3f8gXPlP5LSVAox1cSppQW1sW81+5grG6NZm26uHECuYefTmNGAWvQJeerFI6h0871MJPAVdt4D5hOBQXuvyyujdLfJ6GrCaz6YhegdEcQaoBYUXQewSjdk2ISTkfrHboCIYBcxRN2WPsrekzZkCOIDks73CNaY2dnrAfltRf7y2JU3UXmtqrusNmzHsNKATMDCKyhXsSvU47BKd/SrezXI7cRPbi1tRhqAtrpEE1KML1KdIxkheaclIYQBdVVOJYUQ1wICjh8tg8yhB0irktwZ0cy9yCfuzht3NEgpi6NzUjQzZrKqPnJLhH67oHCe8NhyRfI3XEGoql+Dl3MeI+5qNADLM9KptqSdi1OhMjRng5pdJodTphlTx+JdFnro+YDnvP+oLY8a/2WJwPUV3eloEIMJmNyaN7ZDbM7S4IgDyQJCbG3U9vxAjMs99IbPRmOWiZmXq9naVRHJk7B+5cgoiWyTS26rGCwfD0i6X7xiHahDDuxSf3MhXFvjt2Y32Km1Ig1HF73DSyCR1LDQxhlGjaYa5p+IVKKtiWGlEbHMba+mUQbqTQ6A25YVoUYG9xNF9osFPY/kfntSBHEzqVHuaUQ8QmzOhHHLpjG2szLIQtGq61ctwYD3Wowp0XygUyyuCUMCy6xY6N2OgJmIYAlTFdq5Ilgc1vJjJK8DWSmpNXV7EVWSFZji8j0i6qKbO06HXaZwOPuSMuF1E9tC5KqvoZbJcR0DMeKV1Sva+0djBWgBvAvocsDC2tNoDJlrXZdnzHlUsug7QnAQTXdnJBObcPJzGQNprgNq/BjOruaOHBsrfaWa3X9U5RpevDDjSFv9hudTEyIdZThlLCRXrgOTeEPCtYjKYLneYINl1WYtFsm5P26EezBOh69DgGrBBUBdj8t46w0AJWAu7RgmVtJ3hLLCKaLfwqK9PER8MUMy2LdWJshio7uVokoa0vD8lqDEOckCrNZZQxDeQbEGYtroCPFAguuu8dGrGaMBiwLxfQ2IWE/UKNLHxPyVKXUii6z9dJ0J9do0lLF0AAysLWmTlt16w4NDC8IDhtYOgghYjvMOCVubQlRFjllQqsS9v6C5fB7bVXFNixfZlITy6b06Fc8wVod3/JT293/IAbHsxK3UNVekUsUnUXWDq7zY6FoOpXmGGEtjZNw2RwkupJVacMWUDZaAN1iNSI1RuPaN43OyeYOq6qkBWl6wewALZlyqNQ8HFe8VkScv2jSOuSNpNV2JWr1sPLK/8AAFqGbekcsiYnWB043JaHwFo2DuGejiDcqJqxatzlJav8nxGxplrQAhJEThRboHioMfl9bL/I21Ppq/YyzV/guaXgG0RklXKtmHFp7o/suAQiLC6Z3lO8oxo1desLBZmCsxL404Cgx2IZtwJDshsJ8wQrbdWzVN1mxc9akKx9xNamXO7VV7GUAyXQgCPAt6MevUcSximyDBfDKE4+IUblRZ+I2ZUe6ArpLNsaun4l2D8sXCW0dRYLE3I+BQL3PokMxYq0GFEJCzTtEGPkmJyNIobe0GBFdjEUNd1zO3Sa7niqOHg3SMJNFCqaHiOamEDTVAaI3GqWqt3o1cugKrSvxCUOOh/k/wAM/wAlqIaUUGM3dbBBzHULR0iBWn4ILr5HRixrtS0i4U2plTit2LhC9K1EeYIxqHEeNSzSe+H3YEVAUBCpa+1zY5jSmooh1qAoQCnphKeJohO0zYmGu6Jvjn+RcC9er7oavMOi8oiNaOvMaUvZA0Rp1hnqzNuwB3lhBBqz2UEWcgawMbsy5Zs2L04gTCP03mzHv/qWLBfrmPU8pI8g0uKO6zqvA2vSyb4Ui+2+RtCMAbDokoZcuI1gURAK5ivA7cSqlXoHIIBIbQtUDSV0bNTpGwE2KXI3NKB6/wCpTGm7YPe4NllQF0abqJvvVDlZutyHQAsyvUOXqcabSp8qE0+j/oQta2uxghplDG0SsAu1hxCKKEbn5g4xn0AShYxzvKz+aoC6TXvrBKtBCd6jFR6SHXkOSOioFg9846kuyHSFG5xD4+ruJf0S5R5ZKHYdoUXDgaezfuT/ALf+Q+pIWIys5b3bsc9z4hSwBoJKMhN9RSyvAbscRdiKi6jQ6EJXQwNDtA5IYb+hYPMeodoC/uhN6SZ6cWVeIJoEo9do9o3PHaZekYM+/wDCp0J2Sg6pQ4qD2z36OzFMtNtmi2Rii0MdI3A4YFcbOrwBzDfZwnk/A0IGlH1gN1CfdxV7gq/xHFDrBXsqNWO9X+YdZ5k1aDVl7jMehmbXVd15hU6RWJRrEZlWVXqqexyRUvKePKN0eCXdahirs5UvNMjMki9Bq2Nr40rqsvYFdJdpVsVj8y19H3jseZ/qP+h/USdi0qHFdCY5SkvgEqCEGjsXFWx/qEJI9YiWJENnvm1se6oZYLFvZYRkHWJ2bpSVu3hTxowAaf1ED7wylr9zL1q/isAoNlEsQ79I6MU0/L5g8qA5aN13v9QBWgFvaK9AMaF7ghKEUaNU6SCfRRwJb2RYqx1+LhZa7MAM0/BAN3r00W3X8kQUdKuuXY+8MAUDVhYKKKS9AkCUXN0awDvmLHqxtWmbgqhTb/Gaq8cmWOi2AjoEY/1G1+c8JWycO9IdYg6KJbnQFTqZzG3UVvBeWEbUEoAiWtVLOmiBasDd/kZqZV2f5Mu29Q6v5ECWQ5Y+JSl3fR+IvFSMWIqo6FRcsoC0xaBOm8rToDINbPEX5vaFJDJ4uBeHm2EX0nOTmfEPawW5ltV6wSrQKvXaVgZVSxi3OY9aRtY8k2qaKAM3vioRZ+7BkfgiNWt8ExZkcKTn4p7sZXUzjfx5CAZKrlbD3qsnRgIWWtTvW16w3sO7vDb35WpqevHeADgre8nrcIjOANhrDWqInYZnr0uodKdSAS2LyRgX6j/YjV+x/sRhY7ZfETGBfS4eHrRqOr54nGoByatw9oF5au6jXuJYFepEMvRoBDDhfaM/4ECjSpi0jwkDWUxNEkBN13ki5m3h/Zyzsf7DAMwCz5hBolvRo3qRWXBbbBO5K5RU+bcPyNoAIbGxOYc53EFQBVeJeQVHlPkQNYAAKojgipjHWMpBhdPycx4hwNl0a0YhY1sNRFmc6x4jG2bxnUAfmWKHW2TVXERtm+QJQ7Or+7rMd+ptL1ICq6GZY1y6XcXV2lYwFvqtVeZo6mHWo3p7iV9iDqPI7MV36oe0NSKCTCo9qVNu0BC4sUPUmgLzsdB+4ZK2ycSqgubMJP8AqSuTjDsqzTqdYZAu+Mp4TNJ6nZq/Wsf77AHA2PmI/SGOstysoINkrEdYTte8SBZ4BA2PaInBowPaCwEoh53R1hI+wdESiawSkCjEDQvWCggB8Xw35IHKqNiMOsIanJ/OsPGxQVg4/qX1bE1r0lH4vakGbYjQeihU3hzQeSFhdfyhyYuC8fQNXl5ZVLDiY86RQR6Bmge8VKVpQTywfMrbbow0+3cbkHbSZ4cQsr16z8Euhuao6BZasooqEg2C5uS6n9Y8/B/WJc19P7xHPIIJ1csFaFsASrNXFqNY63YOVM34jDLSybOt6tOLjYmAbDxGFHEZWsHS9PeNOAE1rJbnGektCqHRgK/b2mgETCfiBmh5f5FWlTu/yauJyL/IOJSkKJm8Z2PMIxA8OLznYlRoS6BMFaDHy6/Fy1IUVLoKBeLsA4Q7SNn7xQQi2F5z4D3iWUckApu5aEFcF5L3XqxG8wtLdF44PmFmfC/5EaR0X8gAvOk/EXe8QRNUIQzYzLtvIB6UTAeXQpAvEQe+GvLQVK1LGDb5Q6eGeFBRbOjAfsZuUkLdqBbrL6EAkY6wurGHjHMCxUsl6aqis8rX/aLVeBok1QQ0w5M3WYY0DWqvzPbjf2YMfCP6gdYNqs/pDwJGXYxhgE+7W3JtKJmdapy7R2FDW1+gRjF1zPEehKH9gqaWZOkOg2yrGbp0v5Rtu8n5LKCNsRVrgc4T2jFM0DC5MvUhRgutMBku2INjtH3uAZMVu+vmUjX5ZSmXCwnxC9FVdHmo0AUD7AIzF/hIIRG3aYv8t3Qf0mQDJAZBpOebxDFQAaM378+8sexQlXHxE2CO4Sk5eBGvKNoV9zMCXzCzV+ROkL0YB3tP3QSntbRVaxfxRGrGj+kIxJoMBW0ccGI42+gGBlIjbZOpLCQ0ANrU15ICsp7yr9yT4vM5Z0WwBBlYQeRpYcKNbPyQXjIG022N07bSmKLQ3ioj/V/G6XwQcIoD57ykQ1fmEut5sjMF2VAI+8yrzoBuMPmX19JSVOu9YYKZjiPjSWq0OVgdEdyDropL3hDegG0OOp0gI6FFWsFtjmOEXr6m18GkOgVGYIYgGDK/8hud1CrNhnnCGneF6fhOh0d4dSwSM7gjTCfC36g4vephLGisrw94WN/0wPaLUr2lPVCNUb2aEbYe2gRsIAR/kGannS9ccFAQvW6Rt7Q57rVb+pT2Rc3mtFlNccQxCAdMzWQe5LStYepQpGpKbtmFM6P/AAYm22VwjitjpAU2gVsS55Hg1Yk0udfZt1hZq4HZkMfNakcC5ZTY4tUc9XrKA2hTSAbM8biZoKUGqxB9tYnP6QfZsYO1Kbcj2gXk2BzoezbtCzGUC1ovHglJKACjV/k3a7iG88gRJAnc/iUcgPQrlcaEsu2YrerAu1vecXJMNNIisStnHE0uDDw7JKrAoORNDzx0h69hBJoM8AkN5QYyWkc6xKF3ZV26EGI9yVGHOsdIe9OiJLVDEEu6EASdtc2+0RBbqipur91ltNR1Zojl/kchMQgZKSYoy3kbqHHSYYpJbsnxUvRbgU1x21gClZwjA4UKVxfAiygGqiUdm9LSC52wcozoLvdTAQF6K/hEUq8pAlvdFSy/MQI5WHZmGOfkslvlqwWNYi8W9kGKOISGnEIvjiHyqVuxohOmox/hKBxnXV0igxHFVaPiNhoCqMvgDaqVTsJNhl6gaB8waXSyskd/zLIKVcBqob6ass5o3qchKwmhggozG5xiO5NuzB7UMSmSlhfzChTiYi8L7L7RbTmoN/mVbvgQd37Mey3giUWBUVrB3L9opugHR+kpXRkAXg61B3WwjxkDaJRNk0qHaWhVx2QBB0SUVmriNSGiUcYRlOeAaWuvEB8r4iz50il+s/sBMsdj+yhkvt/YOIDiqM/MChAUbE3rkh6leIJLQP1LNusBZ05hoTBzDLqr1lYPXu6YGIqZhnBc7x3wFwtsjMkll02hFjLeYp/aGDXSmkpQ5qVz56wwVH+D0iWEAqupSrjpKUyxmVPWKThLTfugFlmCgnRjTSAjzC3pQWJxNzaYrmjKnTaOMkxlfyDVU3I/iBtjD4rdWR4WWE10VFrFS7AmV0f5MhmJ9LHWE1DIjYw0lntFX0lt0yuWCEbeYWTKND8rUZdK2qF0G3UhMU1fcK4qdZJ10qqDFKy6tovjJYKDgfthBlalc2zB6nSbZo1C6XTVYhqXK6y40ssxbzWN4TFgUN6G70IiAgcC7pwdIAYMzeoXRAvOjvDUI9FtRUXAx/ZUGToOfwmWY2Nvy8szYohrpfQIq9AXKhxh0gWEBQuBgPMEOSaZSHjXSAbscdOiPLtCCLQEriyUnecWUKAYOXiVYo4GwmPisjnqvAGVlz76Pu9IlhGpRZV2ilLxEgIoIUJThxoyx23Y4RsRs39qmygxC6uhFX+BEGnADd3jbDsnNKtolIvHMx/pil3mY4y0SGivSm75izcJ0KuzmwiY8ZbTx9OsvlWzWp7zVA9/7R5n6cxGU99MqhpFYIjd+L+INw1FlnQinW6ZmX3jJ2KuN/kq5QZLUdKBdgVNYlXQJsMTEbkrAaJVv3RDjhplqXdPtj5vxDfLug2lh2YBAm3iur80DPmKmElRPBkLghhNgEkeTuZUHIN4Cy+8wy6x/vBQQjGQI0HBioKAbIKq5l6LbUWXvioaKTUWCsXSXU1cqu3GLm5rc/uFp0hQrMDagFFF6XAt7czWGNbp94AVQcOAnW6yY63pTUTFrwRPXtkW9iJErFqqutQrwTdsr0zpVTWbA3Mgti13+YxQGquYBxULQB3Nq+CyzHCIG0Ooph93gXp5lxVJZnvkHfTeXOm4EWdZTb1yZ8It1G+YHVzMFrPBTZ4mEenQ7fDLzph6E7awwNc8faVAxqtvZmMJ8ohUjGWNt86Q7t9iVO6BaKzFoSMFThf3XpEvrPEoPzf5hr8yu/U2BdKze4ZpVeIT+rloZ8EzFvVXQHeUJZAcDa3MoxgsVMDYybP7MHmYdrjeWh2hTqBarhs0Y6h8rRrc3EvP4IolJNcEi1WfUfoITzwonAsEuZRMRNSigZtlIII3/wBDfvMBC0qnyQQjjK5UvFBF1aSq4/OWTEiWbjN4zkcxwx0bwGKkFIwetzikHxZXmMEiNANwb+IE0r1B6xCcGgjdqOU4eq2ekPlPYThNolNTNZU8zVVXcAdrJ/WNhIVpGoQ3u29TRdYyVcjr1Hc6k6fuhDYGHSI5V0ioINgCCFzDsz9QzPSbJ0bIOS0wPfHW0Nah94A8guAm+yqxULN1HtZQrSLCsQ24WpQEs+Bw/A8HWK7hobDpFHEWL6zs9pwxQzGBV2utXi5phGLpN03b+MxyNuh1NerAWxLoBDxmWbei41iM7w7djWNMbA4ebYkW3UqcALvcvt0sf0DzzDqwWNlThW+RiU9i2HVtYFutrWZVebX7gaPtusKOjz/sNVp4j3DglxoErrELhEaBWrtLLJocvWt7g67/AIhqZnjcOsaHM0vRbNYvyxFqXs58kbqZvJmHBO0/koidaH+TIUnh/IDtIGfiUIUmErW6Mrb2Sonqyg6Vxu+0wmptLFUvhf7Ko9Ay72Ji3XVr0EeSDPw0YgjQpGCsfm5rCQ7a697h06MNOwmZg5t1BoK7WvtNOXvUcljxFA1/IQHfKZK8yp0NEBDOvWOIGHMi5ZkcLYpxRLJFtaO+iIeXOx99CJ371Px0mTDSlWzHotgVaseFgEurWXH14t+TRiYDpW176MrEBBbsVMwB3P8AsIAcYEf2K7vExTQLzCUd1l/mUQKDWHEcWHNoDdYagEpPCzuA09xlGxISodrUFmifwy/zW+l/7M3Xqiy01Gse6xMWHufA4jHIGZt3LiQCIrbch2JmrsJpjGKVTNADUIsxveLu+pj/AMNhACtxR6fYLm+g7NPmMr9KdU0T7xMDJAyBh+IuA8HHDL827ixlq8C/BxGiV/VG8AggZG2trMphTgTUSE7tVDG4dmOxgGvjWs8TW1eh/kSPsiG10ESwV+ompSTFB1slzrlDsHlNkQuBN1GutGCdwqXUZe06sUFNS6XuzAGxmVvWDEe7lVeWAw+1MSninKNRmgU6akskLwe8SBlcy7IKBQG1ri9xAyi17M1AeKtgTIcw8HtNbVkphhmsxTTdNDCiXkVYy2ziVa7TJbL9CLls2lQoYai4HPWVmwYb37QsR8Uq2k4B2uNvGejBrmMOJoBuplXRFcGGNicDclE1W7HUtyXCYMuYJYYYU+8zaRdKscpK6AXOPOxP+P8AxEXBTbVXUbsuA3CrPJpHuAnMPeHPDQavjEZFAJCODGXrNDFHEwoX1jppWYmZQf5AJcpgJlVRUxkRcgeHQR8UXKmO5v2i1astZTuYvnRB4qxBxsioeLEl6X82Sy6lmmBfJvAr9LYWjQdAS/ExaIz3iaTQKhutiWSr1LR1f6neii7yw8ErRGpKHO0LzvDgFHyteekUyqdOd7l3Cy1DmixBwCdUQ7m1Yo8LAh199Ib8wELlzH2OrHIz0yD1DTzNdO6tf8RaWNW/NCWwNLXpBa7FlXoHaNspbiU0/diXKG2tDTWJrA4gK/vVjTSOE/yVCLuf5BcCvVVq3TFGfEIDhKXTY64lY9Gpqg/5HISEIui3dgA6lFQON0KDG7yu7FXdqgj2Am7BLzqHpoHykSjdPjl5Fe8C91wMbs50DV8mEEgMvdz+wZewp/ZTSE+ZHVaXFXEXpW9svVI5FpXimM4y0SA0Ut5g9xgBRKHA0gG0bO8O2oK77H5mY2OjqPyaQoQN01gt6K4lBKE6S1IvCjVGdDMgH7lIMSa0x8wTIq3cAt9LiipDQYmb5pDcT096zxgQpVD5qFvYiZCFVBMvGE9xbLTp1sfVEEaUIpgy6wuWXcWVmmSV2O01yho0upQtzIB8QRpAoF6U7DcBhKjal+0sPLf5htT99Ipbp1YmBpV4cFvDcQcA2DgjM1FYHTLHxM7BzwC6rv8AqF5VYRCi/BKhipXvLrBWyFF6u32hwkrvDokXUiUpzqdz9TEFc/wlTkHVR36XUwXyp5iFh+WZ9DcLERhJak6Cke6bRW0wc+BF9Bw8iJhhNeQm90SKhtxgdP7mtxbhbgs6Es7RTRmJ1PU0luBqPmKKxRax6zP/AFgAWvOsDH3KC/aU9s0OPZaSB6NFKR4TrA6sBnAzwHpAMiEbXK+LnXPDp4l6pVn2byPSASyctOY5ZxF8QRZrAI9gfAeSWRrnHbJeSI0Xdwu53Kr/ADNy7tq9y4q8hkfCdYVpkLjgqN0NJ1HZlsD0FsDo6wBcFiYhaJudOkaOKgjDp2gVoLC6z2njHrNHEai7EBjGjFHnOqLvYmGq2jcgPG56RCmoGDc4wHQgmUgD5Jct34lWZICszRZygd1lp4l5YqDFRFZRz0lyp1YronL1jigvVlWCO3LOuDgOhGsGFahwWxuz7H+zKPif7MdwQGLf+oCo6luMZYOao9AIKIUlyxsq3Xr/AJLDstv8RmmApBbuyhfWBYq7vSpVKkCRkjQHjMPVjibBxexHF5Zl4GIFjuC/mbtdzMnY8iaufQEcLtglfyAf9bbF68F4l+Gs1M6useYJWuSllpdnTa7u8pL18Q1CjdCeVFCPHxMHTXl0Fm/JtNM/gkuaWtNMdCJdXv8A4m16H2QAtdz+RB7Mv5AgJ1RwLikTEKLdMW0eXMOulUAoXQbtNJTsWnDS7go2qjg0D2hG0sdPhidWNjiIypctYwfP4lloWdND5/EMc4bgNtNDGr0h3HgJRjJziIsOxqVtgKejDA3abT/SCgu7n9ZUWQCvoAFoPaHsS+GKFt5YB0EnNjkh1cQ1JzGzLzENgXJhlM0xTclMaEmBCMmdICJXWwYjhW8tMRaY3rkOtQhG8D1KRhtSdxv5iuA4/wCpiO7D0uAjhK1UQkDcJUSBb0ax8ojUmEFrzZQotveiAuEJojLhqQ8sHUy3E4VUgQo3jzNMLEeZSq2xqRKg5muIiBuLRWLtZvZOIwyC/kritskYwddu8OowOBwumtkRU5Q0/UYTsv8AiDbPH/iVFdV/xKQzONAab1sQ8S5fBVVKQc7MlExAHIs5xAPOU86Se8UD5S8CUJYYa8QhLLTytYSMdk0VgO8f26qMlZdyc9cw0EoId9c8+8XDwfVRtL3x/wAQGLfrpK/6n8gebbya/EVUgiEOOpDtdw/B1lRWkh/AOtvcpHARmIsXe5ntpHlzENkrE3hmhEXbJC9aIwC1iFCAgMBDUldHpBgnfl+JUYd6aP5Btrn/AIgglG6CpVLUpxO1T/CdIeYYGXEBavPmnrAJsrTbBdGdZThJ0SXJtF4OIIIEw/esvcGINvMJWkt2gJpTtB3eJhIWoy8P13HgfRlQc7P7BgJmtD8wHD2S7MCWUqid0TReGXqL6qMYqx0TiNi5z4EaHSNc5KC1FPTJyQixbUobq76ZxASWbjrLSgz1gtRK9Mk78adP0grgBoaeIPTFoDxiPMgYdkxRxrUpbYMbgOUwMKRHwyjwEXmi4Wq9IXNNIVS7SgJ1DC2mxeoeYUOD3bctLNusrqWS6m+8XEQlc8EzMxtdPKEVpYKmdisEvWzPrtG6L6cR+WUU1uwYgLl2Msd0/EDC0qWzf8n+zMmnE4UKBc1WvfUvI/AcEYvjKM9UMujQDcJd4nzfYhuE5xWsEnG4LKq2LFhiE9QQB2LiEAuAwfM17zv9nWfL+xKUPb/UERvtBn+4ClEqHavw4jOzhq7sPLofENs1A0FsdiXQAaTaKaYEROtEKPOom917EEg2gmmQ8t3MpKWlUYB7DUzLGIPe7uYch4xTT2v8hJF0p/IyD2hf1LlOhp5ZM1l8R61IKrTSNEs2doDhkV3ojZirrVPwQQIMtO8W7HeKsCzWcQUvdENt3lgdi0UrwhfrFaZZHdoiFXI0ewjiznWAGPq/5jRZ0/8AMt+oPrEp3MEBFISLgtFrdGrcN4IDSX8QCivH0IOrgqBNF8Ze0fLapa+3iIywkxLAmvKt2bS+I0NStcADz+ImbgrPQgh3Uu/BGaoLZuUJekUbu5E4WAyDa4EJEWMmHHO3BFC+XiP6PAF7GDeuZqQos7n9UpivCR5GLV78QUfwgzqHKmntpBGXz0drPNS8wJoDufMHfRBwMwoJSuZeNjFJW49NkhgkiaXNTphisaLlHKsNa0xR/W5M2LI/WY9yjKB/Yjc9BECh4zXaPRAFuzjXzXMEJb10MjuZOzLY0v2ghd9Lj0s0tFdK7fiLUlNopUYh3EsBYoZubl2Pt+4g0cOnQ6rMMlWmlrD4ple6ALT0aRTW7v8A5NUBfL/kq5+/iEUbu/8AkWt1Oo9qhXwj6LsNAL5ghBaTPD+GKOkHa2GI95NSGEGCOLdDKxWxpGmVrEvOJLpuTqviVt0sMAUEsW7kL6zLP3Iswjv/AJDv5H+Qd7nH4hrvZBQ3LIfElXLY1H9wy7rJbNA/mdMKNalE0vUZZdAOjn4GBUxMmCXpSYlmliAC6/qAmWGNPJfl/kGh4BgAqHUBeV1xsxPWUsJ8wovN7f2aVAUWQBbAx8DI2dYGro4Gxhw0VUcjsy1ZiPJ0JvKY67nbMuwO3WPMsZudRup0ZqZGrVcJswgE1JQUnd8QXqr4+WxWWCQqCcjktpELte0drT/IXIlwk7bb533qOIYY+YVM6wJTDLHTMTgN5lHbYz8v/AmWCR7kHF3fAxu2p0nwBWIJkdBg6RwzdrcxvS46KGnvEUjxA6H8Jp3efwhFE4AELzodGxoa9JhZWkOkOutw2QKeukOwodwzjjUd5eEYwlBobrwRxcJ6QiVvFgIBTyV/2Ycxd7EljrTTW8cMbdM3W9g/MzO8hXUwY2ZlgGD4hTC++IAxTvUsMGg5I7U0FhR7w9mKsp/IWEKgaBMhRBi5pubNIAYobYZRyRMQLbN3iHgLI+b3Y66pIvbLVcqMDqx8HFzVcn1sRr49ARmgvFzb/W6yljg+jF8uTo/sU1en+0ZcfDJmCxkl5Xbboe8o8BBVuWr2Lhr8KvQwfMA7DrWmvYzGiOUeoxReSRN3OXIJYwPBAQ8BpfTzcv3h7lv2x3gsBqsqhyvdSZ2tVqXmJKaeyINF7IBh0CjX2lTuM2n8mjCtuerOlCCSfS7Q5QPWRS0Lp2qoo2qXtWr9RUXuw+QNR8ytBwcIc+9vI4efxK13uVA+xcUTAG4wNIJwokgpdGM9QIqMBs+JXHZq/wCIUpvOz4iIENVI2OJRkhllMhpEq1yP+Iqt3LE01veLaMqa3Y+Qhlubrt88S+MBVqAlJZXhfW4n2qArsfMzFZDXKIlt8smkVGtIM27RkAOxrTA6jEm2SciQPtV2GGkcF8nI66ZHxLCw1GFx5z/UENXt/sed7f7HcN+94QcgvWoISlqcAHfQjQZO03cya1AkXVRSawcTwuLlVFaKJDqaEIKq64DoSlAmBahubcdan2YygEVou+dvw9IwJGnD+wIpLw/sKr+P/YLc8f7EHKeP9mkJqB9wtTDhkds5rQSrHUbc0Xf8yhsNyLo9YvQt5gLCyiYqD3K8eHMrDRd8vTpHuW827A7cQ9EsUMBquSNcSiadmbjqJ8Qa/dP9g3Ldb/2UQo6C/mCrLmJcDbZniZO3pUFOR8SzfMray3w4iRGjsUdk+GIWDTTV+TrH0KdE/wBhYGUOkU1Ya4QD5jHu8FqeBcoeJXYyTfYVUPH9TW19Qa5MZi5o2fsgkPNlfEKlqX09rD0gIRHXw8xKIpLZupmiRGkdXwaDrUR3W2HCJEnOLGR4G/fWB2EtWHWtyJU7LzLfWJD9d0oiru5gx6xK3RYaACUnMVNtG9t20IZM2mpMd85i9IxYODqbEQw1ilA4Ox13iNliBla2GitV2P3zDmQOvvKX9pgbNTKLc0Z8DRcl70xsfaw5WtAMNTeJUdrtyxVAUcUYhVmBQAWrQI6usrIOK7PWB7CQ/EzcwP3wBZp07RfTkkdDqjdemzp/a7sdzNaGNbuf5BA3BmdzZ/sfrZswIRhW8n8gxpe38l4YniAgU03tGDJUlo1CDY0ihlYNgwGqxHvIMabr2IdlFuPQPaVGpdZdyw6rdla2piOKA6yhoYdYUkwgNBeGa0vq8QT7gdmrQUiGNekYr1FI2rO0LYx/ekS5+3iMGLrb/IQubVV0Mld+gwwYpw16vdt8wrxx1LzZvR+ZTozzBQLuJnPZAHsyoZixOIxThbhQrmYRoPzBx2rok3d8w1KdPVyeXVgnDQN9d3L8TUnhP9gVyb7/ANhMPcwAQ+C4vd6kMPyaRhqoL5aKdyCmw5CTa2cVW5dqwS2oVbqwQLESmOoXSvVHS5S05nE1KigLer2x7zVCuOED8iHLZB9XwYmRmXGUB16SkNNNItbcOSAAsYKAfLRMPYMgvG0LLh5aGsxBlmbZl1C8QVPMmkyUVOajjM6x3GF2fFt/7QoGxHWJcOFuI0Sa8rt0mGFcoq36RUIxQBMBQWjF4tSG5CtLuCExsNf5Mc7Cs04fzHJwEwLI0VpYxfoC/wDEA4Tv/mC083+YMy+/+Yk4omgqrmz/AJT7xitBqYzPNZji/GpSuBZ0gcB3zM9a4yLLI044BiqNCbKFhJdONT9EgsTnXTuOo2o7X0Wg+2+3/Yk4FLlaRzvnr9nClyxG6k1QjbZkraITOLi5Tlpj4v7hoqxYjdywBpbzVqFvStxgQFPE3H3ioHjqBiQglfvJaQWrVR7BGHpKrMDyYgC1/txLun7F/UV/3J1EikMtU+s1NkfztKqD9n7+GPyuoIGovSysQCgGXoOGaFxAWrw/2PVh4bRjuzseI78aVu5q2uVrWQyQ8jbaIi3ZDwVN/wBJ0l3euyh0b16T+x/1Eq6aN/3K3Dn2CL+Yfu5lwnaDYN2NOj5/UCvyGdVdYu3dkdsKNXSPI7QKCcKYdv7n/Fzky75yxXTmPDNUyhtwbC70Pz0aZptlYnBOVKhXOVrpwcvSZedWWnK/UukUuLXWzGZxQMaHUd3HiOClKMg2KaMKm4qgEIWh5xBTSnQsjHuQBcG6SjAW22WUNBRlNLxESAC1XBGeiYvrELu0hiPLD2V/IGkAINyJ0iLunN36RnG1XZf2MBjnoXB+zUdUw2F/EXmBpwhB3KNtH+yqYrdh/sWu/Zf7NfF6XCidCios7sXbMvbtEma0jv4ga1P2y1IxwwyQbNzYSWIxY9iB1i0LgFd5z8PRik/OargdA2iqZAA40Ve35uam0YBWtEGG/q7yvXxf6jVny/6jw/R5jRZho/spMEOMOwXsNX1cQF4SAjpVzNl5AFp71HGkmFUh9F2BqGjMxPsLI6J4jPBFviCHEqwFU0oYSBjpvnMcC0DBR/ktz8TUW2LyPeW/9btBlP2P1K0W+j+pYBhswpQOFFU7yn5pANP+3EKRyRpNhVZ0lT5LB4lmjSIhplqejGbG26WY906FmLUD8yoSInBU2e9Qt+nzn4RCJZvWXM4m+LLi6vXLMm93kwBDdZ2dTQSFpzLyuEKdNVt2hBpp9gjUbgpRKGFq2RcOpwIP7hu1QDIM15hYK3jVXg7hLx3sXRDT4Yl4jzFwQQ1vPVWYEDOsJMl3KtiqwG0GvMwzD6bx2ONhA+Yt3YG8TYYeQYWbz7cxDpnaH/oRR+1GuPmjojEShMexcPORHhS7dx8wkeWxo06U3M3CcU9k5gNdka53mr72NbSp+UdAaQhzBhGc0C+2Cw5hAR1xS6Un3IQv6tMMx/X1hS/hxG14xXQuxijSXbDDZBVTMXTFMvCMiaDddISkFWV8i6xjDTGJeyWKymsfYVW2b3QK1VcSzYsmg3GH4TVuW4zWdo6szo0eLNozRVKz6xLSHKoeILgpC6odRGZCSiErfr1giAnBs2Y2290sPWUug4YP2Bi1teHp1lUBhN+qFW0HVfMAiCAm/RgSbm0Qq0doHJ7pQkizjkqVckfIuhm/ArHeAlPo9IyEGw/yEgPIaOcQFjjKZsilXHXoA8kI5vJBiJT1ian+PQRjO/5UFpLhOaDA7SO//WL2e0xhIEaz/XWH8Wk6f66xStURs/OAifYA8Dd9pS1iRQ0utOZSq5iqBG0VXev6m7Pb+pZOsjPDMV5x2NWwC69YoBoN+YF5KOICJACUfDg9/HaOGEZP3KUXbE8gwDntBd05M/EFe23s6j04llsuzaCs3baBn2ICMlKwOAIsZV6j+wYH6DrMP0XmfeB7x8FQAZ2CIULhHScDWPQfcjaWrU/QjqhjmCC8wyVw9wsowGm+wJ/2OLILiCWqm87Nuu6Hg0bAXzefuYv6X2i9fJ/Ofvr/AJwT9/2mL992hYnh5mAErS0iHGpcord8tvmadmIUTB7s+JbPbqXdZqgrKyzAJdLUEg7dFxvgro6x3GALZTSo8qhpikyV91hHWealH8D3jdUSCMpZXMsABh6zTghWrEA3juQ0M9GbiCrW1eIZlK6RT02hpVnZvLllqX5ioVCXZRCcon553iVr+GUPmMz6hraFu1SvajLldVhFKoYllgdd3ZcW/Of3DFhXu94Fxrwf3HO2AZzCm7gtxdlaWDMTcghMdG1IkKtMCMfxE0n/ANKqzSvERmglRqkQrgCXAKtIA5ut8UsHMlsPvQRAWHylz0Y0x5WVN4HeMo2kquAwM/uMszXJRsaOLu3iPbSrQqPweDEaEgmwxgt2YDAK1YQ3DXUr/DJ7SrvY51GxmXOC8hORWLmVSltOIFMqsSwGApDu0iDZYFqJGIX9AGjpejzDYuiHJ3q+dfeP0A7f5K19mn8lBR7D+R2h/XSWaB9dJQ/CCpZDGzKa5AOEl6ysPtQrwR12l2PEuyqwXTxNU0CYQU3mOtbqICxpu3PeD4CQzd+kKLgOleJbO10IkdYu4lf8HENJHnd6HvHnwLrIOWpGNpJaLe7MFlhlaDhlA6C66e37g2ACAhGZctDAu3RgFLvIkaNnm5r4luo9oblKBdkzVRVeUKyS0ljj/CUUzpfqMxlWF34mpijFZyQZ29o5lC5g2BXVGRFyv/UDq9LulNgLV2jJIsI1e0Dmq+eZg4mQaHX+I2sOL47dJW9Est1iOZtqJWo+51q7uyon5hErdd7xYl5c6wLqdGZXtA0O1FOILq+swVpwgCiqmRfdiuQ5L2HSUxWJxcx2UniK0vgVbRCo78uzxcRsAReCXRfEowtIa1tmbb9pbD5/5y5a/f8AnN39npB3fk/lDWS/ttCucuUNNswk9MCCHOo8Rx11HT+jKOrqQd41DNwUygRzAvI0IXH6cwPHctAM0X8veM12LDv5/kUuJF1zxtBa3d8A1RlV9X5i9j994QBOv95naMIMWuc0D7w4ggpIfEuuskq2pedJp1pAhp5h0wAwNQjigyYmFEsK02wY4thbVjZyJadCpSRUaa6moPaiGcULp0gOi+IpqhAgxr+mYRv9XjhDERUH8mqBmnlgT/FOShgPLdYYuKKdVXvpKPbKAZqYOIiWqUEtdqjPYLdYI+yLxbSTWFA0QFajZJfXYZdLbQXUJqZoqBRXONKNBCguzviORTtSEDMDwIydUGTltIr0RlRUQAANW+Y9MW9NyjckBkF29pheOxtHS5Y62dXYwbaOqiDkXGr4goXDeX8RNAWCG8a1EwNx41E6Ix/YFcE0ARjJcJJXjpGHbkYsaj0/yPqMP1tFz7viM6fl/Juqez/JSo71Nq9mmUrxtVQpzKcGkZ3p5grBdy5XmDy4i+BckjgXd6tKY2LsCsytY4/hG7+/AOfTGcRzvnmUOp7WTS8+pF32xM4D5/ycP1ukA/J/KYyh9uJT0TKqP1ABPLHQqMbNtnRlmBefKjM3sHsnIzCxFcwk2d8kruy8IaoF6ViduYLL/kWU/oWEqLYzHgQoA16ukJilACJETDIR+CFjKdpHStBUtKzAZlpuIXQurlK2cXKObjTD0gw7jVydTpBShnOst6iFdrw2vf0lVGbIBBLTeZSlsM1o+AB1GPszFoDd6+kco6lBXzHeoGcfMUCY5FA3zUQkqwanWiXdbkyL7zrPefYcp8Mm7uz4mfKx1dpqd58Nmrun1+j6e+ajz6S0u80EdfM+Q/E1po8R37ej9dwz6nWfC9P5D8Q1Rm02mqfacJ+k+Z+U0TT3T8s1O0+DPquZ9vyjp6hNU1poZ8d/Efc8k+x4Q0d5odvTU958T0X9TyT4U+D/AAjoTQzZHWNKfEfzNGH5eslpdvR+N/M+Y/LPp+HpH5U+u4ZrJv8AW8fVoGl29V0eJ8JGt3n1fE+51mj6bz880Zo8J9JzPouE/D+59Haa32zPwzUx1O01J8mfPz6Tg9NfCZoz5E1o1To7Z9lzPr+HpbQ7Q/c1+81dk+x3m+flfifWczV+uWa/f9zS7zUzZDR49D9rzPmJ9tzNPiaI0E0e2GjPnPzNPxPyT6Tifl/maM/HPiJ8onxH4mtPweoj4c1nb9x0/wDEp//Z" }, {"x": -545,"y": 460,"w": 1114,"h": 1146, "type": "color", "background_color": "rgba(255,255,255,0.919014)", "border-radius": 0 }, {"x": -512,"y": 342,"w": 1083,"h": 776,"type":"text","text": "","text-data": "{title}","font": "roboto","color": "#000000","font-size": 28, "font-style":"regular", "justification": 0 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAIAAABGuDosAAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nMy9ecxtS1Yfttaqqj2c6Rvu+O59/br7db8mQAARiTikcYwdOzaiDYgIwmg3cmKjOLFDCLENjlpO5EwGoQiIIyA2QlYI2Ca2EbYCkSGJlQSSYMzUDd39ptvvzvebz7CHqpU/at57n/se3R3bW+9995w9VK1atYbfWrVqH/yHv3MKycHM2VcAA4wABIiI7iozEfZsb0YCMMCAOH583LJthJkZCAEZGBgAp2+eaMTfjf42BmKwnQOzAaDJTg2zHQ4AI6K/GkaJAMhJr1MEMAAa18jwnsAcd9LRyAwABhkAAT398eb0GJwMlA/OMIBrbnRp3Ej4mt7sqMv7z1oDY78hIACFcSEiAbtLiPZMyh600uCGnYyYQ6+IAECR9YNR2K+ICMwICGDc3MQpYwDgpFsEhNEYB/ej69a2z5M8sWfQSxYAIDIAyMAynmQxgPAjsw0jABEigkLotW8LwDBj0qcbGTvNQSfTyRjsg575QaTguQdCNipE5MAu20ImeYGinKVRJ9+mu8Fh2yavb9MUemUFCP1wGLs7w2x5yslt+3QmMNUZF9cFD+6EXBoGeuIHYDmIsFdR7fnkC7O9HclNWWhwLGFOd/2ok/Ppd06v2AGORJYhfWJMom81HeRwsPEKxgfe7h4GRkAvtgAA0sqL1dpJJQmto+8FESUAI2twDwMzAXi9BwBgZEj6QQAEjNbEC26ise6f/IbpY6DDllWcNmj9hjHoXAoiGnZGwXMCMh67SQIwidHK+YAAjIDo/ZRJ7hn7XkRAQOZsjAQ5bxHB8ORY90phaOu5R/DV+UlgRGBw3nvcPlpTmAzYfTIYLV0gjJnt7DtTN5bF9DNC1vj+0YETJ0RmmLjDaixaYq2V9JLtns7Mij0XVSBnUUqGf5AJnZdmZulnmb1QJDqa2DAM1oWBkAOyCgPwOuCsiHDuAZI7PMNH8CBILjNgMPfoWkMENtZ2ujFk/tSNm4MnAm/EMUNcQ+cDHLQqsvI5ziE0ElVi0pRM2m9m9t5uBAA8BYTRRkG0VuBd9z7ZSpUhQz4eqyBE7BB4E41Uwp6AoPw5C2HY+T10UCCRP+9kgAfiPrazI6ndMxzPpv13Zn150xbvTxwCADB56cKRug0Fyc9WyiaPsjwEGLgRR1BkECCyQhQEjZ7qKQoPJDMVApjEPFu9H4gLQDSyHAhl77mtdkzLJfnxm/G1METfYEKtteNOS3Hgu59z7BeICeFwgwXrfuKd3tdYYsIUBmxtTSOG2MYRPGVYR4GBY/UeGIXOAGXALNjJZEKZEDBB0L6jOC7vL71b2XOMrdt4CBZ/jvU/bcR2PIyCYDgj4EUGgINs7Osdvft005B0SlnHwIjgRuFYwGStkB+cRBTkY/TRgNExf0xHouIACEAAxHlYHSgl/x8CIiOw/Zz3MjVOh2wmLzKDGeDvMGHOiXGkEoOEZe3n4xnPXE5homyBJwbABEyCXjbRNxhF1RLgSQqtU+INMO86tf3OQHFugyLOBQCDwAkJnHDDOlhPZG6bvRZFmQsdQM6x8TRNxFqhEec43xGAnDyZnkUAQiZkgoj8M1YwOBAROzSJ94hjkYOHncewBs9HKLYtgYCEBMDMAlEAav+wk5XEukAOuJNbIHbkHOYwuI4khofdv+yHz6nJhlToI8KGZPQW4mCM6pMo2Uuybzyd6SSODAAoDG2ft2Fmm/ozwD5iifGSG7r3aGPQPHT9yad4KU03hGdN5hAgOgoEZkSIEcOw9ZHYIRKDgejZkhtCpOZYNKR56vOEyXckBJFEGj0OI6Ua8Cr97LU2EYupB4MXing+Rimj+znXkHTiCSCkJhz/bfgNgAAGwXgY5H2ZuxEgU8GkS/evT18EDiFPIcshxRBGH0xmuD21cJzcGfjE6A10enC8hpBoj4X1Q1yRNgvx1thUtO5RdOwAKUvgeBudjBq9/ptk2nwgh64ZYOO0yut0vDeT1NTeQbQslp4RF0aHHyzmJiDYncCJCWHd22Cm9k5kmN0gGBitCXu7pgaHZw4PaH3eI4ke2b5Dcm/YLAMiSEzivAR9hltto/6vh7UOe7pk7duPCr2cRavubDMjomCXjgg9jxUGERMDGOmzXmsQxSK43LRhDl4lndRAlQEGTuwqBr+Z059o/mBQEERqNEPkfNoA+DEET20pCigLAMmLDfooBcBreDIR4cNUZMJRTdEzNaVgwpxbGcE0d+RMl/Pzw7EFAvKZ2geBskecvY+u28s5eylzMzvZKQDQACEAImBYxtl3cLIgEewLhjAwWY2JdzLIYKWiIE5EnEgWe9rv5LRqbE4m+OJzvmPHEmzzSHL3D9Ty1fMm/zfzJPY7BfWIcprJeoiJs07CE+56CkwmhCWF8ulf/8jEfCMwsl2NRcSIlSk4Gw8W2aHzIVPQk+coTu0Uc8jpD4STR+rh+e9ma4CLCADRRHeRCNCYCenww0mbxvN3WGvCANk99p9IJQBydOl2gkxyc2Yj/JizKHHPmixE28RhyAME64THwyUZ5DM1h04yktZtnMcIxAAAhlGPKHDcCe7CB3+BP/tkK+q1s+vgnaEVEsrCkmT8wTsmkDjhRRgLOGNqfJASOeIV2I1xStkRETwo8tHUlEtJEE4yha5uYPCI5bCIjw7iKvZTyIwuHkg7SxAg+IsZ0KDEIkRbHS4lKBTZmeTYXNoFD7VzYGtH9Eyt4gdVDhTlMwXJVEI+A8G+BEuKXmfiCkRC26DZ7FKUxQyIhgxe+mywphKRnN/nwKIgEsFGAQMjB5uUiZKf+sRF5kPFpD/wA4bREWSInH5mFEEukdlMJInRvY7ZuhQ30GkfFRTANuTmka3xIk9hAgYRQrLIsDfRnmJ/E2MikcN4MZetQElipNmSbYbnU5doMZmTdWYN6LCD9T/eJlhASuDz2pGshAOBtKgA6P8kcPZtY4+U2gxQucff9mlgZPLJzjQWjytZuVhlmukITyxi2m8UXrsSGi30EBCyW1OHKMbepMbwBQEACFmBjTwMIZsomQN7FmLczIQM/BGlq9sDj5zEQmGsk8vOUdoin9A+5rHhEEHZLgjZDGUj5WAAZt7/Omakw8RsWOhSfKkZ9ygHHEbyrmFA/PgYAJUB/ehdQtRhCIjLwFAgsvnmBBlMukHOF7L8g9HMZ/52uhFOI1tIV05yaYkQg4ckeaMY6DAASMESpo7HZjyStLUl2HLdsQqRgSmOPDH8ToynWM0uUSWT+oNIOgnwEbATDUWEwMawEkiIrWZCYOOyATByr+jyYBFhRScTZnkkptPO0TdkBX6gSNnw0PhGo5pzDlAirrP0DKEzApsQvKHrLjIUBmEJJldcU26VD6OKe6CXOHYv1Z5LvnwgxTCQCmI6BECLvPwiFwAgsy833KN7mF+YCAsB2EEOd0sQ7hQ2w1QjQayd9ka0EMxctNOT9ES4i8B2ocynghKVn7QarjFHXgjbMtCLIYBFH58lvY9YkUBl6QlIKgC96gEDABEYgQzMRIDChRmSQGs2QdhSYqMEDe33gCCfLY6UpeYkFZfA4KgkCeeGID52YmA8M/421xQA2FA05tbC7ZlvTAfynDSLs+ZpdVOmGJ4VUXGjaQv3TwRUccqCU0uP6eKulOAJXBc8IcOwPW9dPeFDt4YYdBIBOMEEKWBI282H4G9Ft1AHGMXO2a8RIsoQaWLR4g02K5C4k5QkRkjUODyf+7T41z2Y1Pb6tGRurLxlcn7CP08IhIj57ZB4MB/XZkIAflbACTqHgpIc6o2C4FzcGGBgXLL58+YiEyM/6KxZv+ATgtexoCWUMAQAOenBRnZoYKcDCYiD3FNS/YsAPITPiEjM2mIJv0g87UVzGgZR9dAv+UrKTGNSEfdxSWaPczF11TrOBwaVcoZzCNj2pJgwGDs//0hR7AKOSlgC8fNIf8Lo/VDssDIdHpuhwWerRmA1BGMvDD5qx7Q9AAI0BgBQkqs6sezwcME+wj6FH9cHEvOPkeZk9JZ8Zy9SR5N58NRLcGiHOeIU61gS+GulIRt55AsGaMP+fDRyDhEmshU/eM3jdHL2H5PcT8/ENJ1VvWBzRm0TAiC7gtBRF2PJS305OhCYNMwQIHjSAkYr4WHPGFn5M1a2XR0cBbHxi3+ToGgw/tFA8yDWqyymEur/4UhbzByNWBylOcIEj132YQHHK2RkkNYTJPqAAD5P79Uo1WdtWFgMBExoi2HDODH7x32MfiaOZ8SRKCjBnwxtVbQVIT0Tcqn2MRPwmxf9yCWHif20xT8ZbZZpSATM4wrI4H+ZmYERRXrejSe3uIOrg+6GQWp2Nc45J+Pdp5VDLmWDAkx9RYptKQjbRMOZwZ4aY8rCRF7BJ86jqYrEJFqB0TZN5YgZBvcHmjz2wIAQ008Jj2wTg5bjAt3YZkXy/SFxxBr2yxpD+tBjRGebUXjBi1bWSSk5J2u3UuWrVIlQR51JFtzHFA2PFL+lhp+iCqTVWbbTUKQNA1gRAKH/C34DWCQjl13bcIyex7H7QJ58d46wzCWmnHFy5m/mzOgPODDo155EtytmwvZ7rXPD8ThuAEWNbSQE7G5F1c9mZs1dWmJM3TBQHA8z1z0Yw1scfZjoxf9J58lOXxhmVIs95mN8sF9Qt+5GUpLMspchXdrzHoJt3grBMGi0+3LZYACgQebssrABcGDdKfBA2nLqMhjjBeWdHAE52M+BCGYHhtIYIj7lxS90NJlwRA84YbTsHoQtDT+djplxvOM6RbY226vQnumP+oOe9tENgw/hcGYCAFJH6j1SjuZx0GAqQ3b0GJQ1bhUNSduBXxqPd4Lg5NLeQXFY7d6vHFlw5c9gblKcO8mnbp9WTDTuSRzX9nqfFYwZgglKyUwIAEQIJBAMa+ej06XXQBgD0Jj7I0g5NMCchSsAdv1kQkjTZjCFleh9CbLPZ0Vshjbwd2VA7IebGL3cQnPUvoQIBw/clFCQp2B+ADJBTFDJIEqPR7A1kWkpo/IbvTWL5W0QdQGs8oZ0sqNhj9BxXnzgb7Y9MXDmKCIcdXwdzW9+eADJiEyMe4mIRELM/L6zw0NURERAXzPu1osSJUl4QYBmyg5jViYDCCjDGNI7wKtgEkMAAAsASVAIFHZPjebGpImXTA2YOa+m8djfqhmjmTQm4QFm8Nvf0wupXqUmf6IRAHD7DC1xEWSgqw1CBnBLUT7Qx0RSPSV+/x9iWNsGL44exnt7DelfJ2aYjDQ6hryuB0Po6CSb07mAoAAQnrfxIXs58FNGWe1MMLH23yjK7BnhhpOAMAgmNPP3aSQYB5y1P/01jjrZrRFGDaNjUiAnj8QcJfWnjGCn1b1UAACAbFqZWeBwU9KgX0w/+LqsZAgjKpnBLhkTsiAU5LtkNllV7HQLzJxpQbJkG9fW/DEw28xMqaR6Qp+T3xycT2FAUojhfaJfk7L6aEN5Hrqw6EstzTAIS9htHR4gRCuGuXZ7WUQXi9EwvPY6hz4A8CUiLnHI04MNBsU96G3q9J0ZQ+zWEWsdonJmz2Tf2MOZMViekGYcPD2+M5Fwj0Iy9UhuDg4VARiJnb5xeA+I3wWUUO3dI4AvHHJnIcmwpyN1TImkyTBGL8o00GDLDkQmRAIEQONRPsS6/L0FUYjDNZ1B2+l4IqmsU4Q20Wb+1NDKBe5kLXh2Jzuhk0WUDK55uDIQl4B6E1yWmNgU8OzjhnetHuTnShK0egDn8o5yV+KHkfeLPhsZ/PkI6yZJ8ygXwa57u5B7ekpN3lhPUk/n1sV9PISDO+MkOqoosaUTXghDM+kRbOh0xfGwkcHGvvifT9J4n+1vYOk78hrlq0oZ2OcCI6LVzDY5JQjsJllC1gzogF2cDPDewsoSe+wdBILBsEEvkEOZAAtBOL5yII3I0+zQPi0anRnYzgnPHTqKpmvYpruNGGNpShZHjWP6oYf0je99KkaKDkOEbfowUKQ4qmh73RhSlxtmfRAKBkuReOfEUjiiI/np973gB+3705Kn4gs1Qj9JbW+g3vecWD//KS5VBfoDoAJAtziRcm98pDYi1KL66tih9iajQekZnYuho9dVPkaz4WvEjAEiIwmFAY0QJpHZag64AimHKTDkxx289WAjZUSqJOBUJMQuNLBb45G4hpKsVPSzubvw7VuJiJaM3WxOZGOZU4HMKB2oaBapT5bDDI980NmV0Zodh6kK3gaTRnyEsUdIkNEt5SYAB8N4Ar8d71LHC14MXL8Dg51QGLexZ5qWHv5a4KafC3/NT50bbxCQ56Lrcc5gEgoyc24qouaM72cOPgTGVhWd+bF1RhiK0jEYHwaQRK3R4AcX2nbxcUKI/Wi8cbQqDbbs0nseSvjJEIozAe1z3jimYxyKoKc6jCjCqtyN2DMm4jwKl529Cch8wA4/wAQUZIYYrbMdHanQZDY0cV+QzHEG1l2noT7PGx9IgUEw8wPH662bY+pIJ50jd49jCEwYAmjMXeXQlcWxR29mEAgh8yipZKZ1aP6TyeYIY3oaGNwGyHS2vSmggDTyY6zDXswiwZzEXcPhIDCDjELpLT0hZjst3ByhAQBmAiBEArB53t4YBHZFtRP2YshKJ6mx8SjxHOxY3Hrl0ZdlThCHWHg/AWwmjqy+N3Iqct+PHhJ76QybM2OYuOnQrNPU4Kwia5MzLrABYACRF9G4vWJBJSEQxd54e2p9AJ6rYvAIGQSCKO7JmBG8bHicmz/ilQGD7u8zxhQe8DpNmSzuiy6nj1ATMchrRdsXVGOfd3zHxyQ4dKg7G2OYC5SD5wNN48ZtZolceGF5biVpgvA0OE6JS5yJM1AAJn06t2+ZJYTU3sDgJGYGOCkK9uMKPjQOx/cC6MqAbROJ/WYYDS0zpQEnmPzyIE7wyZZkDpzaDDIFUTST7E3YGhZwyHD4yVCGOMQjtZCJCYbetx0cdR7oD9oJn8n3F+hI4A2ABeJx0JOSFGkDNIM3eYyF2G1oe0fqNjzG4fvwqx9FeCK9LUdZSROTAI4CNHFJUhS2OF6z4dHdkcVDKbPte8zmIZs7T2NOBHOHid4NOgvyFPAJJBIc7IOPJxDSabQJPns+n5x9AGOQPACXtbZibKsbcWhWAUNJTJiEJHqB1Lkxc8AC1lcQgtPi6LTSltydY1uV+1jOVSu6I8CEu4PwaWJZJp7J0/HRAjr+eAFMYF9YxORwDvMss4WRHjUE+wLPKdgZDDaHV6n/nyq4RiSiICODY2JNffw1eGX3mnUGRc4+SFsfz5EdMZ7zVjNNQ8FA4LyM+vNWCNxMpQbW/8tBENPC+SRQnzD7roVogCMMiGGGlwDNI1ZkFobTK2DrcaKvSM18fMiCQTsmRzQnwNSxJTYae/MFZQOrHKQyy/NOZ5ec8E/IU/rgpHr4vZOQGpUBc9xhIg/GQCAAVocbxr7GlkJ5TxmyEX6RJPVKIxY5DsZPo7FPcWUAHbPBhUuIKCdDHD/UgbI6PMwhULRvZBw9lulK5kwszfGZIVxGhzziPXlQHgLBYItylLJnJF4+xzFZYnWQnbCHlwYEFQ3mDCAxdex3R0DU6jCoAd/HjpHJh1kckFAmoPFvULoog/Faol5TXBjkdgaxBIZ2UoUJrQZqU9/l3muVUhFITRO54Upm+CcPSviXgmRLNCT8SQ/vtNhpHQ+Efnx/pmD5EKLttooRnpKIyMYQ+d99wGCeU9sfuWQQgLk3iMCCHMcCi+IMJS4rCjEbv3xIabkkJJNH7vc2AOxbh9DWQYYXKYy5kLogSDTIDyO7K0r3JBMpmW3fWjbj4EqdQhXwyGg5L/s8gQjtEaJ/AwSEvfshYLPn8+gAQ6yddZrI06DjSdiZXgoAwXuqqB5BdYNhAjCAlDrJeGXc71T6K57JPwec5QBpzFVMtQzg5sWv1DnnQxOU5M9mMz9AyymRllfMLNEtCPq0ijUDmKJIS44Bn85iAM1AAMggCKWBdlCLx8kGPz/mbO78XnD/mK88BwRg4ZYtLcusCBnvL6ZY4F0Vx+88mqOIFgIzBtKUYGX3yknjDJWLcq1XYQA0fv/+1DEo3EitQDiTmPOojGEIAdybBPygUxszrHuYpmLocMb0pF8pGJUBwB4YIxAJV59TDpe9InXQlzMuvr4jQSHoAeFw+vxnCx3cFp2Bo8uG6t1imiSEOOPO1qUx8th22EOOMlEMGF785xvyvBpwwlo+W6+lA0cGN0YD77FmAm9cijdYwGSrhqcL2SW+2Jc8YAouE8XIvGbixXBIOTiSkhAjxUVJTXVmyfweE89ApztpGVQIN9wDwOz27oa3O8QpCY6II0RLCGXE+HsjznYlhWYe9XBuCNjnGsfpltj3ZFgy6VfTRjBSHrJZfhYi/nK4MQPTOc+tFFjdwD1aFMeYgMr9EcFwgPlhrZnVrgSuZhrFSBMVjZj8OkKyhQggRREhLHDwGsFATFEzsyBbNTlUtdGwnTmGhOMuBhhsMkl7B8CQgI/bcvKcRs4bBv9OKNd8RFwDnMZR6sP5fLbsdduXL6tOdSDw2S3GhcH6+DqgAPLAksPiDAdgwQG4TCJpC4yDdYhyaRnIqexipkLRfHJqSseiNpEVTVxVUlGdmLCES84eRc4MFzcCeQBscTTtEfe30QJ/jF5Mmhg5SM1QOAXBrk1RtfeQqVymd3vMyibrzJFk3Fy7N2cJZCbsXdI3GqqMjqSXGHMneUO373WqODnm+xDYQQ8KisS5anrzHySHk4U9TrUJvV2yuRxEv90jgfXoZNqdT9x/8FFRvdGqCoZKqrjyGqqH0LUKkMpsIH44W9bocrCgic8MnMn5nEiz53DqUrIYZ3+/wUcFTnAIYe2HzLlBtLCeqmw+wgymXyfH62crfXoA9vK2/SSnNouTM5nxfTt9GAcqe9dDgl6QE98MDlmLxsAmSjT7HETm3we5lDFfEnEE706yGyLi9AuOPpkGVgSdiYco31nIEeyIT03lk7s/JIxk2EKMIFMmf0NLJhDoFIndg16HyJPNTvjIMTkDWKGoEsFXCodWwVflBK/FVh8SD5xl0jFsrgpjQf91nFuysjFwxlG6wkAcOYmWp7bPubsgM4hh8R4BkrRtAigS3g3UAxKNGYL3EYjIBgNxQsdPDaQrEg8IbMgy14u1TB9On4nNjfgYfBYiEoIgYEaJwOQhhDPgI3c8oixv2k2/X5/mxMqnFtG9H9Ug2O0xXlzZx36eUIe0Ag3BpSSfAjcdiAnJ3xjkoX+Lu2UduA8Qc72h1+BXEMGXcxt09tiKiK8E4/EMRo44WnKowsApN2IdSngk3u7x26S95DDAoEXgXZ+zhIOa/IEi57V/3lS7DGigOgUdgYGQWvQJx5WdGQr6lP1HyKQcctGaQI/TX11iKOnYCaDMdNFxLdwyAkWOJeAbRUIga74RhK8J1w7RJ/sgvWzl3Y2shSOPvfRGNJUOyepo2DwIGfRk47GNTY2m/gcc5AIvo1GjAgUJpo8Ol2gEwHyfVo/QP5gNCgEAxEC9fezhb0m0ejiWqMOIOXJJhIw5SPYA/wSVjiNMO/JcYj+/CG7HJaKv0PVMSzaiZfLNvlkfgqcKn2zuxex+dz1o+NDQ5B1lEXLa+H5NCzcEZBibze/yLcDAFZF345Ij6e8siZ80bjM57MYPktxWNTs/nJRshbk3U5EoDOCBv539pcn4dTDs1OeGDv2gBzzCZM55yLT0zokeI6WY/HXN7m0pfzI+hYHvIxPLHAEMjGd52j+jDeecbni8lmefIbhnBzijqKUKuYcPKQ6wz6TuOn0ALQIPNHBQJOfwfD7muZGB58XzXcH4mNANK+dDWJT6w1GbiBJzV4x59X9QxDEoAkBmMAaQWJJ98RYwg2HQejJzCABMDl5w8ElBAULv7jP4YGc40qE/nYQEBgCZ7TblFKYHuJyUxCYOPJnjCLMS7jkXlGDjpOvYWtJARrBtQiCyYQh7ASDJOyehnm0SEe2OUwgb23LEkXPHOpSI3FPDmBU4uX+9QdljgwYQ1+OxaMU8zVMaaJWQfJgYXaUnC/falL3gPGXx/iM60sznewPA2T3Pa8fvwo2voIiw3oOiQZfpwQzG/7oruWp+CKEbBx+aWnf0w2QACDZkD62IwIx+WwMEdx/+H2E2/9X+IHdQiWFMCF54GCDUFE0HcM4QBxGwd7IH6xaADZ2DD1cS1JYWCIVtjMDMDqOnr97wfs3lRB30zSxAzrGEdATwC5sOwmHUrQBshuOFqYnOzYrdSZEvdMRUuOVVojcJXPfdgQffkVOR7Fym90HxGCbuP5LRZUI1fuZtHRF4DUn0NRigkcQOSI8ggxnJrisgIfS+gUDgnkGGlKm7ZxBsxDtdU5a0KOleboYGlePOuyBoXjM5mfVIhJ02ThFXZsMyWYFgBDDMVDIbnisjEbQ0ewbbwYa3Z1kiKGiG08oQkXuD7zk+eonMcNkXvQkCv9ln/AOGuX+AaB6H4AT8Ap8fQ1SQwPRM1iH4VfQt+KYDi+KjUwo5FLac5sHNQx5nH7KVGUfISC8moxrb+1S2d6B6eStDUXZrN/Z3X92apSRmBsOoDZtRQiWVNgBGBkbyXycQlLs5qFs6fgZ0uDLs6pmwheRkKm5aHBADkXHR2wQ0NXBAmOKnxM9iQvNz3Dd5RDUADKnsoLe0dvT2lQDe03nsF2J8tr+O4TRARyQZhdq/BcSOEABsiGCiuAc6GJL9cOx/Nc7n9KeCgUD5GNsE3RgCUNfXBLsGMY+vEce09N3j6ohvQ0iT8OZ5kCxF5gM140y9cUJDAnGDWZ4Cvi6DwX68jG6xE4mBcbdfUqKXQCflBjLpHSHg6QYAIIkoXBMDFBHC8rjTBBhGNjUVSu9NAW2CbpS5HrRvv46hwmAUCODdQ2JoEy65R9DTY9d74n6AKGWArrLBB1XumRhoZTAsooKsvC/RSeemslKjCcZP6v+eoMhOb0wFRI4996m82WCeMDkz2LHm/P/AdkE+x+lcDLOjo3yxtUoASbZ37KhC0NYAACAASURBVNfefa1elALe7pjW0YT2T/P49J+cbuyz2t7bH79y76rp/Xu5MqmyRpEBwTAbZm2g1bDr9bY3TW80QympklQKkISFAEEkgl/znMW47zy6n7S6epjCGlkNSK8l0HSAQoLfHUDZ9EOOUhy7XV1fbp7zdiG9hF78vVcL1Tk2rAoJd86fHvYS6A87zAdYzkFcW0KBkZagvkkUx9PvXAyO952EMrHpd3Dy7Y/Aw0/z+eljiK7+fz7Yr1GkToIBjIFOQ2v0tuPemKvW9Mza6N6gIDTGKBKdNp2Gs20rSHSaa4mdMfNClIRVIUsBpSBCIJqYHwwbP9jWRU8QBslj5AM1n+YaMh3RF5eO/GeehIx/0w+DKDGjYdRRGMI4eGA7JH89RJvDDT8Mw8R4TnDaJDrPasPh6PUJrBd3fu55u3Df+cH75fkzFc1/yqL92TnsEgEbNp2GTpttZ3a9aTVfNFogdgYMm1LgrtfzUm07ninRGiMAAVAzS+RW81yA1qYTghkvdloSNVe7UmGnTSFFLQiRKylqhaWgQhClwfjbbevORTo5PwqdB9G1RTLjiAuTv/bTWN/SKHyCJA8WkzDNk8ExeZFejEoSd2JOjAjcMwh+rxUC2mQ7gt2EZFXCuB97ZtJoBDBO1mUljf7ujn2B0e9OyMd3py1+BtryWWoGJgdqoUb4zAyfONk9umoUiUYbACil3HVdIURvTKd5pmjd9nWhOm3TELxr+3mpDLDWxgjShtsepaT1rltWsu0YQBeC1o2eFaLpzK7rpRDPtloSsjGaoZJUKSyJykJUAktJREAemgEkWSgGcsvozwsqIOqQc4IuT+UASAwxMK6pP+8Yh3OJ4+BoaUNt9EgDhw9OoKQEZ+ZQLKYVXAhnI2Bgt0WKOUBEjDGNHEfkn96Ro+zP7Jh8fiCWnxnNn7a2JO8V4vAsB7jMcYKuWsNA67ZXkgjxqmlnSvRs2t4sSrlptSAhEK6avlSKge3KpjZGMwBQJVXTd5WSiLjtTCnEZdNVCpUUF7u+LiQzbZquVKrtDQMXgra92fYg0PTrDgCUQAImhrqQs4JKgbUkJVCRsFVC4HRkXD4HI2Tl43jPvrB8hj5Gfn4aI12r9X8dDETH1thI4rRw0FqciKxyO+0XEiWxjo4GCwDpKrlPzAD4DAkGV4wI9s3WllHs5zkh7NM8PgtK8rbHZw99BR/8nCO4CPaFM4majG+1/3LT60qK3vDOmLmSreG2N4tCdhpabZaV6jR2xszA/+gIAwJqZgYWiD0bA1BKcdE0SFQpedV081JVhVi3XSVFIcWm7ZQQkmjT9YJIEW17TYSKRNNrYkRB620PGxaCELDvu0JSKcVCiVlJMykKiZKQ/LqQlQQvJNGoQ8wHOsAOXimmDdpUUUz0CXEXC1iX4fVkEPDwSDWGUC227NaW3O/Pst/OwLZqISS7nGlzKj9IYAwORJSDAbqEZGDXPz/HcwId+Iy0JXs0RUpeMVwaGhPz8c66K6TYdkYQ1IoabXZdv6qkZnO26Y5mlTF8tWuqQmmA3tjXuLJB6LUxhhnA9LqXRiAWUm6ablaoqpIX292iLmul1ru2UKJSsul003OlhGFet12pJCJtu04gCYmd7rVhJUVn2GithOgZm6Y/b7TYIAJ3mhF4rsSilDNFdSFqAVKQICJgvzkyKXsNwgdDyUr8hkEPlSziT1c0k8UC74smikT2HoOUmk+AsRN792bK0D6A/WGtNFOHmQJPZvmCk5ReJkJOL6TWY8LhMzfWnz2L/9w+4J12w6nIe/Rgkt1/E83w6MNzD4F0tWvrQhSErYZd2x9UpQFzse3npQQAZGi1mSMww67rQwlZ76o7oSyKXdvPyqIUcr3bFFIQYaXUxbo5qMt5VVzt2s7omVKd4ctdMy/LeaG2Xd9zP1OKmbdNJ4gqJdtea22UEozYdT0DSCnYcGcYEYjEpjdXbQOIkggRul4XkmYS5oValnJeiEKgJKS8dsbjE899b51pFG+H7xir8nHsZPYdVo32ltYiAHB8KYZbS82A1PCJPd0l1UbWtaH061YmVnBjvDUf3vDzP+MDpz7v1xNO/rALG5hjFPFp+sz0wfTzxbapC6kIGs3rXXM8rwzArtEGjBISAM537ayQgABgdm17MJvZSem1ttBACjpb7+pCGeBVXZ6um8N5KZCkoNNts6qLWakud+1F18xn5bwsr3adEDgvldB8uWukEHWhOm3ON00hRKFUr03Tt1IIJbDXutNGClRIndZaG0ECEZveMAMStgabnXm2bdg0hSICkAQAelEWq0IuSpoVUpLdnBADehvg8JBDAOHtcE6nMt2YzJ1GZ8X+vRkhXgA7eW7DnkdQsbxwvOzzTjK0qV4FBJbmshgdvLQt5gEQTH9OefDP8uDso1eTGFczg4E0gBgeKYaC/DPsV4OJzw7fwrIqzndm0/VX2+baYqYBeq1PN7vbqxkzaDDrdjerlvZXipo+lvfa4mhENsAd615rSQRIALxuurKQUtKm7c43u0Vd1YW8avpnl9vDeTWv1LZtn15sD2bFvCy3XXtytZ1Xal6qpjdnm22pZF2ortcX264QolBCG7Pe9YBcKskMbdszQ6kEMnZtz8xSkhTUaWZmQiAUm65/S7dsTCGFFFAKrCStKrkoZS2pUFg452DXK0z8cQQAyLHNQGQJIe6bAQZfG+rX+31+yVbQOGfENlnr9SKTzUHaemLSE3Rn1SPsIiKXSOZkn3r2T5SSd3gM/Mw/1SNJMNlPFi/x73LDSxqc5oHqhIFwt2Es/vW8dfcwQqv1xaY5Xs0YGAw+vVhfW82YCBgudrtalY5aZ1rtzglgw3bhCgAWZXm5aw/mNQIczKsHZ5fXiwUiLmfVs/O1EG2l1KJU6x0/OV8fL+tCKURzcrVdVGWhZCHketcBdLOqWIiyafuzZjMrylVdtJo3TYcAdSEZoO2MNqZQQgrRa91rjYCVkgzcGmMMSwFEQmswzAJBKEmEPXPT6XUHp00H3Bo2yCiI5wUtCzkv5aIUtQKFSJRlg6M/cJoA3gmEONB5DvJiG/ZQMzD593Ig8J53EtnW90rixCVnomI4ZGsC9tZlOSl4Z8fzVQLzQPfTOYZuO35npxLDVFww589vNfUAkAh6oDy9lD7l9cFHa8mqlr3U9ubZ5ebW4cJK/9luN6uUEsJapov19oXjQwBAxKbTSgqINs9oZvtrFFWhTq62y7q0rx2ZFcXZ5eZwMQc2x6vZ/dPzG6tlIcWsUkj09Hx9vJpLAYeL2flmt2271byc10XX65OrXV2oSomykNum27RtXRSLsui1WTc9MNSlKEl2vVk3LTGUhUSEnUNfWCppDLedZjZCkJTCaG60AWZBhPbdzcDMKAUy0HlrTredhkYgCkSBUAqsFS0qWpXlvBSFAIWEyAbAiTsYBqb4Hg+0+7vQpwlcPO72Lca9vu7uPSCK93itQfbZzqufaE7lRqZob9D0lFA979ivsM8Jst7Bka5B+DedTFOHmZPe1+VAGVJvAHvUJmAnSPTBli37FVs2DBRUk/nZxfr6am5dzKbt1tv2ztHS9nC168qisLkeZl63bSlETCAi9GzIVyz3uu8MSwICWtXVvScni6oWhIBw82D18OTiheOVQCqVoPns4cnFjcOVQjioq23bPz7dHK1qRXS0qLe77uRqs5zVVaFKUJumW+/aWVXMK2UMbJpWG1NXxbyQmmHX9sBcFqIuVW/Mru3YcKGEEIUxZtdqw6YQQkmh2XS9McwFESliw63RwCyEUEIZYwxjb3THuDXwtOlZt8xgDJeSl5U8KNWiEItKlFIUhIBuoxEACPChd1iziAXgEKYiTn4W9/vb30GY7jsZigv69ZDRA15nPq2F9TE1UycB4Dn23WvnPv8A+9xDxHkT66ADyBS+UthWOaItqkqas4k1FxFlsf0NjSSIvHm4vGwNAGvDj88vX7x+ZG8D5odnly/dPAw6fLndLQ5XLgQ0oBl6rRU5CVlV9dVmd7ioLeS4frB8fH5+6/AAGAjoaDF/6/HJ3RvHSCAIj5eLB09Pbx4eKImFogOqn5xdzstyWZdVIQslLzZbzeZgXleFMEo0u+7iqlvM6rpQzLxtu8uur4uiKiQyt9psdjsiqkpJCF1vtm3LbOpCFlL1Wq/b3mijpCilZOa2M73WhKCkQIC20z1rNKykJILeGGPYMBSEsiDD8GxrHl5t2bAiFASEIJAXhTiYqaNKzUtZSRTuFQHsqpwh+ukQxPu1Q4fZGIObGQpJDDxSU/gcaxrelzW5vvPZOQIoSTagcXrVy7L1DLzfRaQ0vQ1s47yH3GOkX8H+IPV+RzH4CgzOdQCAUy3vgrxqG2aBCAD2PZRvPj29fbBC/5Kxy11blQW6dxMxA3SdISBtC8UZAKnvDRdu4uZ18daz09W8stC4KhQYs2v7shAMoKRYLhb3n53dOj4CBCno1vHBw5PT6weHpSIkvL5cnq036217/WCBCItZ1bT907P1wayqSyXroirVxWarDR/M60qpUqpd1z273FZKzKuykKLTer3tNJtZWcxKYRi6Xq/bnUCsy0Io0Wlz1XTGmFJRVUpjuNXGGAaASpFQotfcdNowW8BGgL0x2hhgqKQQksBwb8CA6Qy0DZ40/SdNA8ySUKKpFC1KcTwrV3UxU0Iiht1AbmuYW6EwYXqdReO4P82XlKBbbWT7up9g+RIxSxXBvpXUPmvjRJNY68/aEYLXWPM69A97j/16wKOvOLo6UAzI45MYUTjikhucK/DKAOCXDqPn9p4nsycm/CATM7B5crGeqUJJCsr29Pzi7vUj2xsD9NpIspDKpRYUkWsaEJAFkdHQG0b/+vGb1w7uPTx98eYxAhDioi67rnt6cXl9tbT7c24fHT98drpazJZ1yYiHs9mmbe8/fXb98LAsqFaqWsmz9fb0anP9YCkFLeczrc3Z1RaYV4t5VRZVCW3XP7taE9Gqqha1MMy7tl/vGiVkXaqqEFqbXdt3WhdSzkqJAI3W611vjCmUrAuBgG2vd10HwEpSJaVmaHttJ72QQgrBrNvWaGBkUyipJGmtNQOiADSkBCDuEM4u+o8/uWBmu/xaF+KgKg5rdVCJWSELARLZ/74N2tfdhIg7Tqur4iXPe4BRABODE7tDy2oIRklkcvm1PfDonR0+aHC5Ge8cgJldFOHl0wGbid1aiWdxpyZUJb04oQnJmUx5OHskPTNwFOS9H3s3i7GOxylDgMQWXpN/2yYDbNr+arN76dY1vy8Jt7tWCkEotOMyNJ1WSrGdKrB94c7o2noUZmSqyuJyvT1aLux2E0VyVsiL9W45q20i9HA5f/jk9OLyarWcW2JuHh88OT03bFazGRLMykLJw8dnF/OqPFzMEHA1r7u+eHJxUQp1sJgR0tGybjp9fnWFSAeLWSlFpWZtq8/WWwRezMpKybJQTdudb3YMvCiLqhAVyLbvrzaNYa6UqgqFYJpOX2x7ZlMoWSkJwK029owSWKqCkHtttl1vDAjkQkoCpY3utDGGBYKUglAaY1pjLIJdzQoiYcAww1qbi4vuzfMGEQSiAK4UVpIWJR3NqoNK1QqVy4JhYGxYI8lEaLwxLv+Av/3gYvCAbwbvHFZ29fedHDFJ4HMO7He+DI9QarpPK962r9jSOzoTWo6OBd0GJJO6EQBwv4ZtdcMpR3iDUag7sNnkoB5OYYwhouCR/uovPfjVT3zqpTsvKCL0PHnj4eM7149LpSxtBvjJ+eWsKBZVCeA2mm6b9mq3vXGw8tzjrtePT87v3jgOWM4AvPbWwzs3bxAJy2tt+K1Hj29cO6pVEVj7+ORMSnntYMUAbAwgnF2ut01z+9oBkUBGBrNumvPLq6PlclaVdh910/Vn63WhxOF8bvcjamOudq3pzXJeK0kI3BvYNW3T9XUp67IgRA3ctLrtNIJZzGpJwABNpztttNZ1oVQhEcBoYxf4BWFVFQpRs+m10QaAWUhRCALgTrPWxprvopCCUGvu2ebCQQqhBDGwZraVnuDjSW201gYBKiUqCctSHdbysFazQpSCEJlsRRnTeINXsNfhA9hIPS2JiWHJ3pf/p1GEy/6YoBL+BicoSVCcGmzv4XyWi915d3KsV3mEMAgSYJ+q+CIzjs/6chv/LEEkMnEUEMLxgJocdPKDpnAbAKTq4Zu6/+T0+tGRJLQvsGLgptNGayWlw8WIyHxxtbn2whzJ/3iGZYAvPCEAZpAC265zlKABAAI+XM4fn5zeOj4GAEBGgjs3r7354NGLt24WStoU861rh49Pzx49fXr92hEhEuDRcl4V8v6Tk2uHB7NSAcCiqmpVPLu4uNhsrh+ulKBSypuHq03TPDo5n1XFYlYRilVda6OvtlutzXJel4Wcz8oZl7u2e3a1lYh1WVaFrAqpDV/tWmNMqURdqFJJZm66/nK9Q4CqLOpSEUKvuW27nWFBpJQoJCJAq03TamYjiMpC2iKXXpum1QAgpVRSIkBvYNf2NrQVJJQgADba9MAChVBCChKIGuDpjh+ud71eI3BBVBKUApaVOpipg0rVSiiBiBgMm6/ZYnQ/NDCVy4IROIMY7vNgMS7chT5c5US10ItlDDc8WLRNpAXVmZ4kZDgXGS09OvcUFCOR1KAbtq3wSoLsZAy13cMWASJ6qO8UxGuC5561YDbwyGKPqB5uGMxcSlHMKvQBIgA/fPLs9o1rEA0QMwD3WiABu99msQmbttchyAEAZiSEy/X6YDH3CBUPV4unJ6dtv5RC2uwHIt2+cf1TDx++dOcOkXvf8rWDg9Pzi/sPH925ectazUqVt46Pn56eXRDevHYEgEKIG4eH2659+OyskuL48ACZ66Ksi2Kzax6dntdFcTCvJeHhvO4Mb9v2fL0pC7WcVXUh60J22mx2zcWmL0o1L8tlXQBDp/urbdvrvlSqLlRRSDbQ9+aya4zRpZRloQhIM3d9v9XGaFMoURcFkdCGu14bZmOMFKIsCkLojdl1vTaGDRSCCqWQoNN622u7oVkKVEoQoGbdahOkYlFWgpCB2cBFbx48a5oHl4RYCpRoaimOFtXRTB3Oi2UpC0FkqwHsQvvH7p8n8ukE0xjWhu8ez+aFsD49BVFORCAicvaoOkrtAESF/dUD75CkgDJvN5B4J7URJ+UnOah50O0s/EhjidwgeJ+AmLdpDNvf6hycpPQ1CADg1SP0ZfvV2vzo//34vOnRJ6h2XffG/YevvPtFdIYKAKHt9b1HT1++ewvQ/XgCI7Sduf/s5N23rnurBsC467p7Dx+/7113/YiYATbb5s37j97z4t3oBhmuNpuT02fvuvOi/xFCRsTz9dXJ6elLL9wlir9ef7Fen11c3Ll5069XgmG+2m5PLy5uXTuuSsXGbea+3GyvtuvVYr6sZ+51EsxXu+Zqu5spdbCchbT3tu02TUuAVqMAkRl2bdt0PQMvZ5WtSWOGru9brdnosigqJS3furZvu56RSynqsiAiYOiMaVvNxiByWRaSEBE6bfpeGwZgUxaFkoKAe8NdrzUzAUtBhUWEDJ1m7aqnoVSCBDFD3/faMAP3vbFioLteSSwllQQHlTqo5cGslMxgAHoD205fbNvTdft0024ave3ha77o9ss3ZmnMHspX7IRETJUa40TQrQ7xSFuCKPFUphVi3BwdS7DF4ekQfmHwCOzgSXwcQuTNCEiJHnBc1sBUDazvCAF3PMkwVg9tjIhux5/UhgQxswlv5AB+/Oz01vVrVl61g3qw3jWllFYLtB2TQQToux78GhYzMBspRNu2mo2wiX6DwFwVqlTq7OJytVx4veGqLKuqvn//wQt3XmBjSBADL+uZQPHGp9548YW7UtoUP6/ms7JQDx4/WS3mB6slEhLDaj6bV9XjszM4N7euHSMhIR4s6tW8ulhvHzw7OZjX87pCgoNZdTCrLnftyfkGiQ+WM4E0r8p5WTa9vtjsDPOslLOqnFVVXTGzWe+ay76VBIt5WZWyBg/Ato0xulKqLFVVSWBoO325bbUxkrgqy1klAdhobvq+McDMpaK6LASgBu56vW1azSwQSilnUjBzZ0zTaA2AwIKwkEIgAmCn+85o0GDASCkkCVDUa22MYSkBuAcwiJsd3LtsdL+RP//bT68afblrDRGSKJUohDAkqAAhRYAY6WElOZFVSKx2sjKQ+4Fo3YMCBOXjqEJpX3FlBD1S8fKKIXSONDl7GVvwJwGS3252oXbQjWQUAMYYRKcIgXjDDIl6BH+bqkeInoxx3tmAexkhA3S9Pj2/vHntmtGsEdq+J0Ip6HK9XdSV5qhJViO6rreUeI4gAFdleXJ2cXxwkFgXvHPz5sdefXVWOytuLx0dHj19+uTBo4fXr98U9s2nDFVR3Lxx+/V79168+6JSCt3bwMTtmzdOzk7P37q8c/sFIkQGQrp1dLRrm/tPnszr2dFyYd8YuJzPZlV1fnV1en51dLCaVQqQ6qKYFcWu656cXhrWNw4OlJRK0OFibhiutpuzkwtFcLxaAfOsrLCipmvPr3Zam0LJ1axWSpYFGTZNp8/XO6O5LuWsLMpCMoDW3LTtlW6RcVapWaEIwQQVYmDTL2fVXBUAYBi6vm+a1hhA4FlZ1oKAuTem7U3PDMYQYa2UlMjAnTZtb2wKQACXSgkhbOTTG0OSUKD4/X/8O1VRllWplCxISikkUaXkTKkP3KwPKpHiokHAkgYhA0CCowfSOHsysA74hyNsQ7/AE3q0L5y3pXA4bNne688HNUhNP9slwlHJgPcSw59GshI/9B4M2mgiMWIIM7MQBAC/fO9y2wEzsuGnJyezqlrMakuiJBREwPjg8ZMbx0dIgg0yINi3hhl4dnF57WCJ2asOsSiKR48fHx8eOtfohgzGmKvLy+ViniyIYV3Xp6enhFhVJYN7IZ+QVM9mDx7cL8pCCbu9FBBxVtdC0KNHD2VRCCFsDlIKOZ/Nd03z7PSksIAHABDLopjV1cXV+uziSkopiRBRCDEvi1IWp5dXF+u1VEoKEgSVUou6RMCLzW7bdohCEArCqiirsuy1vtpst7sWAYmEJKqkKJVsuv5q12x2LQAWUpSFqApVKGq7ftP22643DEpRqWSthFKyabtN2+263jBLIUolSikkUdu1u7bbdL0xXChRSyqUEIR91zdat73WxiglSykKKQRR0+u21602zKaQoi5lrYRsDAujBWJFghQRm9Zw03UbwE4bTl9ByZlKhL888AC+NCCkgwbuYqAYidRFp0MD1WLns1JABSEqim2EGpBBIy5bYJfPx78PZowN02F03iCObwdtzFg9gMEYI0iEIRABABvGJyfPPu+VDwjhojebJ2GErmstVgb/A5YEZIi16TxCdSkOw1Ao1bat0ZoEoXs/KyPCzRvXP/6JT7ZdVyhlTYsV8Rfu3HnjjTeQcLFYgn8La6nKF+++6/79tw5Wq+Vq5VEo19Xs9u3y4eOHZVFcP74O4Cpbl4vFbFY/Oz1DhGtHR0oIBGDEw4MVa/Ps/MKY7vjwqCoKZhCCrh2stOGzq6sz3c9m9aKeCYC6LGZl0Rteb7dX266QalHXgmBWFnWhGOBq215stkrKRV0KgUWhClAAsGvb9XYLAIVSi7osy7JCZoNd311uWmOYEOu6qIvCFkF2vV43LRjDCKWUpSpKBADotN40nTW9UoiyEBIRENhw1+qGjTEMiIWiQhIRGgNd328bw4Diq//Ed0lBmnnb6U6bnTaaQQpZCfE5N2YH1fCNcn7RHt745Me0WtSFzM6HCAEAAM4evv43f+pv6vraC9cPg6BD7kk89Mdue/4zf/snX328e/97X3Qi54NoxIEuWUnYcz6kYpPzJp7P5Nr4AGPsDYxhIUbq4bzH6AEAbdXJe5tfeuNy02nDcHJ2TkCr5dJ6GJsMNAxd15+eX1w7PjSMFsiB3cRi4P6Tp9eODgHRuEG5F/uut1vDUNc1+gjMutqirN+8d295eMgh+wdk5fvNN99cLJdSKSKysRyRWK5WJ2enTdfN5zPLEyIiQcvlouv7p0+fzhcLQSSIhCBBtJzPpRQnp2cEsJjXpaRCUFnIw+V8OavPL6/OLy6rqlRSCiIpxbwsF7N503VnV1dd281nFRFJQXVZLOoZIFxtd5ttUyhZKKlIzqpyWVdFIdqu2zW91npWFZKoKopZVZZFwcybpts2LQLXhVLWwJeFINq13a7pNm2npCiVqgtZFqpQUhtu2m7XG637qlCzUpVKlIUExF2nm163XQcAVSkLpYpCCkFam7Zne0lJUReqkEJetR0jS8RlVdife2itYvVsN09H9A3ADOfPHv7c3/vbf/2v//f/6Jd/7d/7vr/xn//pf4sZjO4/+Vu/8ltvbb7qj3y5F33+h3/rR/7Un/nzF7vuff/qN/5vP/PDptk8PTm7fut2IdyvSnzsl/7Bd3zkR/7GT//ktZl67df+0Ye/5Vt/5/7pRr7rjdf/8UEpYvCAUedCyD6Q3KAbAw14TpANIWaYSE8xA4uRT2EGs0c9jDEAWS8GDLPRjJ966/7nfs7nhLQ1s7EFXWeX66Is+x5s6B68MgPoru96g5KM97n24RvXrr/14P7Rwco4ZOn0oaoqqeTp+dlysWL7g082gBTyxXe9+9VXP/ne97+iiABRa2PXmG/cuPX06ZN79+7duv0CIqLRdt7m82VRlp/61L3V4cFisYrRG4rj42vn52dPXnv9+Oh4VtaAbN3karHstX745InzM9Kth9aqqFVxtdu9fv+hILp2eCiICFEgHcxmxpiLy/W211UhD2YzIQgBCqlKhV3fPzq9MMxVUcyqigCUFFIKZmia5t76lBnmVTkvC0FUlwUC9MZcrLe9YQSsS1WXqpRUSoGAvdZn6w0zInBZqKqQs1IhAIPpen25aWyJYyFFoWRFSGDjnG69azUDzQs5l4pQXDbtyXp3tm7appeEc+/+GcAAGIZ7ZKjYwQAAIABJREFUr33yO7/9W7/4X/y87/6v/urn/yu//8aqfOU9rzy89+pP/LUf+Oo/9GVf8ns++Bf+ix9wkmy6n/jB//Rb/vRHPvwd/8ntVfkVX/kH//e//5N/+INf/Mp73/Pf/dQv2Kzib/0fP/u1X/sNv/Hmk0LSP/nFv/OVH/ra9335N335F7/8+77ijzx99dd/+9W3yL3pyb8H2joaBCK39hJ0wEXSNj7J4xAbclhPkCqPYTaGraxjZgTAGIMAgghyLfDqIUYBTBZ+hENJKaS8vLw4WC0KJSUJKYQQQikpBSkhLi4vD5crpYSUUgmphLQ3kBA2RyKFUCQKIZUUSpIUYl7XXd8TkT2jJBVSlIIKKd/70ktPHj0kQiXILjlLQZKoqqoX7tx9643XmJCQlBSCyAYDN2/elEo+uH8PEZBcZR4gVGV196WXtpvd40cPAFkSSZJCCCQ8PDi4df3W+cXloyePrBe3cySlfOHmzWuHx09Pzh4/eaZ77V6YgLCoq1vXry/ni8cnp4+fnTRdx8yGDRCulvObhwdSiMenZ4+eneyaxkJEJcS11fLGwZIQTy8uTi8um7ZDAEFQ19WN1eLGatX3+unl+unZxXq7M2ykwIP57Hi5OJjPuk4/Prt88Oz87HLdaS0ErWb1albO67rvzfnV7uRyc7Hedh0rIed1sajUrCw7bc7Xu5Pz9bOL9abphJBVqWZVIZ+utwwoCAuiupDEDEiaebPZddqbKgAA+JVf/+gbF+r7f+x/+gO/9/c8+NW//6M/+CO/8BP/5fd8yz+Qh7e/+Y9/2+bk4Rd9xR9FhrNHr3/3d3z7T/zsr/zQT/zds//rR1971v30D/3Fv/KJ137fV3394hMP3vf+9wKYX/zpH/kT3/5dTy833/onv/n/+Xs/+uF/5zv/zT/7vd/wL5d/8Id/4+VXmi/90v/2G7/r+37gL357mhILEC6khNOkVn7aZUjRxxD5JXb1VNkKeFAbM3QRfsVfayMEQdgFFxQUQGtNQgwy2tumW2+7N954433v/5zNrrNnfWYQDevTs7Mb12+2bR8p9Jrf9XrX9MgCkh/fcV7ImGdn5weLpe8IfQRHB4vVpz711q1bL2BSHgEIVT2v68Wbr71+++67QlUBABhtlgfHV5fnn/id337Xe98nhGDDAGgIAPna9Zubq4vXPvn67bt3qqqyv+zODCDErZu3umb31v3788Xi6PAQ0f4cLElV3L5xs+u6x89OkOjmtWMil7Euy+KF8nqnu5PzC933x4eHVVkiIBEu62pRVcaYs6v1ydV6VlZHyzkhAtKyrlZ1aZgvN7uLbYPMR6ulkkSAR8uZDS4vd83TyzUwz8pyWddScrGsAWrD0HTd+XqrDQvC1bxWkpbz0gpC2/ebrjONYeaqLOqyWM5Kmy7qtG47fbVrbKgiD2czl2FnbLXedNqwERbt2dDST9+HPvSVH/rQh6zJ/fmf/butad58av7a3/nFf/2DX9yevf5FP/i9f+7f+LKf/R9+6M9/z186fOWD/+uv/OoXvv/Oj/3mT73/X/j8r/umP/bN3/T1P//D3/Pw7I9+8AOH//Wf+5Pf/2M/82e/+yM/+D1/4Td+/sf+1g+8+h9/34//h9/2tb/xC//je15+5Q985dd9+Nu+7Qs/8G4OmSuI25RCLG7XN8TAAdhL7v0dlBDvwl5jGDx88nKCQdlcnJ15FLfJwBgjxAS4AgStNY1TYAxS0G63ravZrC5dGsg1yQDQGmJtytIWPbjNpP46F0IAG6XIbQxFtBE/M7/rXS996q17R6uDoGxg837IL7700q/9k1/lW7eEUAAgEBlYa5ZCXr/1woO33jw7eXrtxk30LhglAXNx7YYqyk+99smXXn6flIUtRCBEJJivVkU9u3/vzcPD1eHRdTteRDTAqNQLd++enZzcu/epGzeuV1UZ0plSyls3b2x2u3v3H87r4vj42OZuDIAQ8sbRsWbz9OSU+5OD1aqua98qHS6XDLzZbu89elJIsVwsSqWsRtdVWZdla/Sjk1MwXJVyuVgKQgBWSpVKGYD1tjm5fCoJ6qpc1DUBCCEWtTTIXa8fn14wsxI0r6uqUIBYFdKK1G7XXa63AlEKUVeFlFQqWSgJwNow/uWff73tdM/GMAiiqpAEaN8o9jWff/2lozKXB3f8v7/4M/eaow/9oQ8KQmD46P/y41/69d/xhR948dX7F3/mu/+zf//f/sZa+U1zLrmlv+ZL7j5bftHu/ke7w/d9/w/+0O/9wrsf+c7/4Fxc+/Cf+ne/5PNeTkQriyg4C0N87B7FLTusAoxSs+5Bu0w++UP39gVVNE5mAUTvMVwWss0aZiaaeEP+X/nFe//nP/61l9/7clXNgH2NmPeCm+323uuvfeBzPtflsIKnQAA2H//Ex2/dvH10cODT3+4XjK0P+fXf/LUv+PwvIPc73rZFA4CG4eT06ZMnT156z/sAwRoCv1SFPff3Pvnxo5u3lssDABSOSWiM0cY0ze7+m6++9PIrhSrTSk0GNMacPn202+5euHNXSP+TTIgILJGM1g8e3FdK3bn9AgmB4R0LAMx8dXlxdnmlpLp2fCyECNlIA8zGnJ6eNb2e1dXhaiVsZ8SIBAy7trncbLUx86pazeeU/C4EA292u8tNg8CzqlzMawGuMKfTTARX292u7Rh4Vhar+Yy8FTUMndFXm22vDQLUZbGsa0F+Cx1y2/Fu19jXBpRKzqtKEOBf+rnXKimlsPwwhpEZ1m3X9vobvvjW+67VAFkC1//xFgMBAB9+7Jf+o4987wf+pS/78Lf9sbs3DiEUd6C3cMw//t985H/+5df+tT/81d/4dV+1qgtIFktCyyYs+WUr2s4CsVsXz9dlrNiElFTebljFAwAaaY5b+NNTKx6ubacekwrJzFprIWRyEQOP/vLPfeJXP/rbn/+5X0DkpMZvkgPN/Ojpk2azeddL745hk72DAZg/8fpri8Xy9o0bvqLO9ubSuL/10Y/evXP3YLXy7UJIcBvDv/lbv3n7xRfLskZmpYTVHGZmYK31xz/2G+95+ZWqnnsI5rwrMzfN7t6rn3jXe18uqllGFbNB2F2tHz546/adu6qoCikRfNYcAQEuLi7OTk5u3by5Wq2cajEwMDIY4PPzi2dPny0Ws+PjazabYdMVCPj/8fXeYXIk151guPSZ5X11te9Go+EGwGC853DIoT9RK/JESpQo6SSdvMTVcknqxJV2KX06ne54kqgVtTSiGR79cEgOx3tgYAa20WiD9ra6y/uqzIyI/SOyCj2GVx8+fEBVZFZmVrx4v/d7v/eCc16tN6qNmibJkWAQIcy9/Xi9+6o3mo1Wi2AUCgaIp5gCon6dcl5rtlrtDobQb+kCtjHAoKegA9Vms9XuQM58pmHpqpiRXChNOG+2Oh3bAZyrCrEMgwhICyEEgHLWbjst2wEAwL97fr1HPrYd6nAGONAlSZbwBw6GB4Pq66dil35901Tb6zHewCaBPZ++5RLOu/u3/rwz8566ZM9K3juzF1f8vDOLmo2f+ymDez5+XSwBhAHgt/QeAABK3TcH7r3Xx7/wMzPWr2l61zF5LlGsWAuLc6FwLBgKYAB6+3QJ8+acrWysESKnE0kBFL3aOS7AGK+Uijv5nbGRCQFA994O4KDRrC8szo/uO4SgIJG5J7SjlGBiO6216zOD+w5IkgK6HL1nl5y71F1fnIsm+03L4nu8mtBrMEY315ZkWY0n0wh5Mk/PbjnAAOTzO45jxxIJIsmcA0opghAjxDlngNcrlUqlYvp8/oDfC/DFXSOAAGi1O6VyVZJIMOCTCBF6MOpSWSYIItuxC5UKgMBvGLqui8ciKAfOGWM8X666jBOCfIauSkTsmQUBF99ertcbHQcjpKmST9MEccM9r4xs1603mxxAjLGpy7LIt0MAAUAQkrbjth2XA0gQNDSZIMg45N0ukt3FqRsQw+6+4q+fweDnTG7Q/bTXC+bGwd21XxyLX5/5u+EZAIAAdomlvaoqzzlACLFXlfHWruP1FFMvngGMcc7fkPjr3QPv+oc3GIB3B4LX6pFnez7qDeAEw4Bp9txal871iK9mozY8NKIS8rpn4n05MnWzY9sSwTciMN5LzKJQKJTNbsoSwtBrbrgXi0qyP+DzN+vlUDjCvZYg4mckDABJMQdGx9cXZ8YP3EQw2vO7cQC4wsno5MH1xXkE3UAoupckQBBBSAZH95XzO2uLswMjY7KsYgghwr1LS6fTjm1nd7YlWYnFYjKRPSsFAACghMOhUKhUKu5uZ/1+v9/v71oJBABIpuSzjE7bLhSLCIJQMKhpGpCwmDc6UTVFZhxUqvXdfIFgHA76xQxFCGEI4pEg4LzZcUrVOgdAlXHQssRPjyEM+cwg55zBUqO5XSwTCE1F0Q0NYYQAlLBkKH5RnlBrtDgDEHFdUXRVhoATglDE1CBEHmkJAeLA5rzabNkuA6KWaM/E7M3+Pbm5Ny6ie80G9QyDv862eim8Gwfx133KOYcQ4b14as8YxhgAe8Xqr1v/+VuyUr0xEFDGQDd+2Htc7x+UUrHx05sWBHF6zhgnBL3ptnjv8FTfUNt1AQBdkOrdL+OAMdZotRiAwo93d46+QWgxDmuNeqvjembFvQwp67abcCgrVqqGbkIAoKjUBl56BHCQSvdfuXROUg2EiHdGwGC39oEouj+cWLh2uX/8AAIEiAQm54iI3hEwnhndWLnebDajsQz3alUg51SskpovBGV1YXY6FEv5g2GEIUGYUtblFVE4mqpUStfn5sLRmOXz7VlrAQNcNSxFN4v5Qj6XC4fDumF68ZCIEREKh8OMsZ3dHGM0GArpus5Zt7AZAk1TVU1p2fba5hZnPBAIqKoqHqxIcQYsk3PeaLWXNncAEPjKFP4XQajLsqZI1OWNVqtQqUEATFM3NU30WIEA+XUNAEg5rzXqpUqdAw4/98yqWKcpZzZlrY7DKAUcGIb2oZtiQ0Fl78TpTYc3xMqvi6T5Hg/6phfzKjFu2MaNAPXGGf7/9mER6byfE3KL1d2LOt7ycAAAZRRBCOHPG+CZx1syV8IWXdclZE9T8DeaIacu/YdXspUW4wB43TIBBIBBCBnnLduevzZ15Kbje9tDeXvzcQ4ArDWbG5sb+8cnIGAQAq8zutdiGwIA8vlcrVoZGhmBvNu6H3it6RjnDIDs9malXu3vH77RWAoCzmCz0TA0jUOwu7niOjQ9NIoRxBA6ros96hIACBhj2Y1lCFC0r9971CKuACJg4y4D2Y1lRmk6MyhLstfCxyNSvKvd2d6ilMbiCUlW8A3n7VXGcEZ3slnK3Gg4qhmG+A4P9QEobiSX23Vs2zQtv9/fizHFdOWcc8DyhWLHdhRFCfr9MsEYQSG5dznnnFMGSpVKp92RCLYsw9BUEWwib9tU7nJYrdfb7Q7G2FIVQ1cxRgh0+VPOGYf4Pb/5CUp5q+PaDoUQ+HUtaGg+TVEkNBHV/JoEelwp8ERNEAl7F/cCRbS412l4mbjuy5vZ3KM00Vt/vjcn+PrPu6O6xoMQgm8eAfa4ju4JurZ641u8yPv1A278uWEe6C0+Fefooi+09/3eHwAAZwwidHqtbruikyeAXtNBr3dapVwEEIWDIZGUESorKDJsCIrIKpfLxWMxCPZeG+rdiawqq6tLiURfl19AvRsV12EY1ubKkhUIypLMAXBsB2MMIVBkSdyYbvlLuW3H7himTzxTb1sNCAFgCELTH2o26sWdTV8gJIiMXigogI3PH8QQba8uyapKZAUhgAUSAYBRhiGyfD5ZUbc21my7o+s6QgiICgQEEQQQIsvn0wwjnytUq2VZlgkhYgHugUNDN03TbDabudyu3bEVVe2anwf/dV23TINxViiWavUmxBAixDhAwGs3oyqKbhiEkFK5WirX2u0OIVK3mwgEgKuyZOqqLMmNVidfrtXqTUoZQJhzTjlgHJBsuSFhbGgy6bbUoiLaFwoi5iUNUQ9Jd62l+88346U3AA8vnNhzhtd9zvdE23vqWN+Amnoa2y6sukGteQcwxgQq7UIjvucbxCGMMYZwDzvt1Zx740RyA0L4etC3514YBV3/yd80gne/BhPStmmz4wAgVjwvDOcQcMa3s9lAKFrvOF1f60l4vQWSA9tmjXqlZTsezQehWNi5l/iGDAKn097J5Uzd7K6tQsTl7e7HOY8k0rNTF8YP3QIRdCjvtDrYK8cSFwUi6ZG1ucsM4kAoCruHespQCAEAZiBKKZu5cr5/7CBCpPvr3Aj6sGZE+obWV67Lhi+ZymDoSb844y6gEEIAcSI9UC0X5menI/EUllRFkjHqpmshgBBFEwnHsbPbW7ZLk8mUoirYgwAQQIAADAUCAb+v2aivr61iTGKxmCTLN6YRhLqqGqrmUlqpVHL5gqHp0XBQIghDIHhGHSv+ZIxxbtudfKFoc6Crqt9nEIwRBAgimYBw0BcCgDLWaLR2ckWEUcDUfYZOLF0BnDsus6Horg1dl9ZbHdtxWx0LQOWtcwQ9pwF+DtzpjeEAop8LaFjXNogg79+CNeJvFXB7r57BiVKNnwecOAeMM8A5IeRNR+8ZQ10s3NPPOYnwUYRIb6QV9pyuF/8oMtKoyEl1HxEHnAPKaa1SHBsb1xQCujtBd0nxbryPAEFYkSWRZ0EAAAhZt7UXgpBz1t8/XMhvJvYf6YmSu6pewa5zQ++rlnZbjUogFJZkwrv6R8/XM845Hz1888LVC5FwSDd0CDy+E/R4fM79vpFoJLK4MNM/Mqkp+t5bFrckEWl44qb8zkZuYyUzPKzKahcldbe8AcBv6al0enNtrVEtJlIZTdOEFxFXyzmXCTYGh6nrbG9vqaqaTiQUWfbMEQHEAUcwYOnJWKzVbK9vbSFCQsGgputAxG+cAwBljGOxKOe80WxuZXOaKkeCfkOVu3kHCCDQVSlgGRyASq2eyxcBgKapW6aGkdjRDsoIKz4j6DNdlzUajc16Hr/7Nz4hYSQTBAGqtzqVRhMwHrb0VNA6kDD9GnkDGurSSwC/CU11x8BeXu/NiGsP6OKMA4SEY0S92EU04IFdMopzjhDqgbq3OI8XdWBP+vA6vNOd+oxCCBHG3dXzjcM4F9TtW5uHFyABTqlLMHnzkrDX8XUJYvDqar3pMO+n6c47xrlL6cbq4sDQOLohrOecgx6lwTljnG9ub6USKVEJAyBgQDQz49y7HqgaxtL8TCI9BEXO3YMAnHPAvGcILH9oZupcMJrmXl//XltCIA5CCFmB0PXpS4FwAmHicVfCQwLAOIQQSLLiCwRX5q4qhiXJknASqIu4MAIcAtMXQBJZW7wuK7KsGLyXmO/ePoLIFwjqurG5utSsN1TL9ECngOUQQggRwgF/QJaV7exOvVnXNBUiTAFgXSoVQiDJJBwKqJpWKOTyxQIiUFNU0pMtQ44RUhXZtAyJkN1CqViuMMYVRYEQMOb1KIAQ6IoSDvhMU2u3mrl8uV5vEIQwxgACyDiEQMJIk2VL14jLaKNlV9s2ZyziM2N+nQBIAXDFqtslf3i32APBvdKe12ER7gEqjiDEwlRA97A9L8Y4AxzfQEyvg0ze34wzvpeMetNZ9rgOL1B64wjvv13ghF7Hhe0ZAABwXdezUi6IpdfvjccFtqZivfe67r3Oc3jPQnTcEVdSrlTztTZzHUy85siMM5fSWqXgtGu72Q0MkUimuq7NqEMUQ8Brypjdbua3FpdDfklSutXysN2qISJ7eQzAGeP1wtbMlVP+YBxDzCDkADDGOq2KZgQQQMLSEOfTZ57yhZKSHuCMKYrMGXNb9Y7T1KwIQohzTiT58smnzEBI1y1JMz27ZaBZzmLDJ6sGgtAIhOYundZlye60gqlBQiSPKGewVNj0hVOEEM3wzU1djsVT1fIukXA4OYQg4pwjDjrNSrmcj8YHdMOq5LPNWlFGeDu7EYzGfYEwhBBDyAEo76whxQyGY3a9Nr21FgjH81urpUK2b+ygpZuAc44QcN3VlblQMqNr5vrstUogCDhfXZ53qTs4OmEqujA3t13f3N6OJNM7pXxlR1VVrVmvzS/MGpYv0zegEAQ5oJTmc9vljhOJxMo7634rwBjd2dpaXV+MD45k0hlNUbB56L7F9fXNbLZVKTVaza2dwtbOztrW1mtXLh5JB1Ihn5DBiuWcMSpiBsY4Y5xR5rguZZR3ZX9coCIq3mGccyr2C3ccfiP5zcXEvXEg54xz13Vdx/GmI2diVrmu69mP+FLOHMehlPacuEA+1LVht/2ueMexO9yrf/Lsh1JKXWfvMEpdx7YBBwhjzxI4p64jyDSxKgDOqetQ18YI762xcp1O7+QAAM6BY7c5o4TIwmpent/Z2c2eefwbg/sOywQTBBCntUrxzOPf0AgZnjikK7KmyLJMitvLW0uzA6MTmiIpiiwRlFuZXZt5LeAPDQ6OWKZh6qqhKktXzhAMBoaG/YZhGoamKfnNpZnzr4xMHIrG45bf9JmGpqoXn3m0b2Qslkj4fIbPNMPR2MzZZ7c3Fo7ffk86GQsHA+FQQNOU6dPPHDx2IpVIREPBeDIRCkfOPvuDRqNy+Ngt0UgkHAoGQ37qtleund935FgsFo2EQ5mhEcjpxTPPIxkfOnwsHo9GIuFgKNiplwo7a/sOHEgm4pmhgWAoVC8Xz51+gUh4dN9YLBIKBX3BcKheyZcrueHR0cGR4XRfXyQRb9ntmdmrgbBvfHxfPB6NRMOReHx3a63dro9PjI2MjoTDwVgi1ei0Fpau+wLW0MhwKhYJR8PRRDy7vY4JOnDwwEAmHYvFkpn+fLm0vLqg+7ShocG+dDyejCfTqWa7JelqOpXIpOLJVCwzMFTvdNZ2sliV+wf6B/rTA0ODiUTcZSwQCiZT8cGBvtGx4aF9++q1+vrOFkcQf/j3P5UIByaH+g6ODfUno0G/WaxVC4ViLBx654n9UZ+GuzgJQUgIESU1IhMkih5lIok3xYTBCIlBYgIxRjkHEpHEsQgiscpihAkhqPsOpRQCIMkSwQRhhBESeIMQodcWOIW5roMgkmQZYUFZIWERkiQh7y0IOHddB2MsyYo3CEHOGWes946gjFzHwZiI6iKBsBhjHHBJknuEGGOMUhdjiUgSvDGMQggJIcLzQAhFKzNCJIS9B3Yx21lcWTSj/WPj44auqaqiKFqlUlzO5g8evSPTP6CqqqKpiqpWG+1weiQZiymqrKiKJKstly3miv0DY/39/ZKiSJIsKzLyReqtTl9fHyEEEwIxwZq5sLqmG3r/0IhEiESIKitKMLq2ND80vI9gQgjBkqxZwdnpK5S2+wb3CXm9pCi6PzR9/lT/6H6JEISRLGuR9MDUhZPVSql/eB/GBCFo+kK6bl0++2K6f1SSZYSA4Q+nBseunHtlbXWhb2BIVhQEUSiWNC3f5Qtn/cGgYZgYoXA8OTA8Nn3x7LWpc9F42jR9BONwPBXwB69cvug6TjAYJJjE44mRkfHlxeuXLp/3+QJBn1+R5XRmwDJ9l65crFQroWBY05S+VGZkZHR9ffXMuTMuhpFg0DKMgUy/pZvzC4u7xYJpGn7TGB4YHB0ez2Z3T50+tZXf0Q0zEggmY+GQ31+sVle2t9u2Ewn4h9LJsaEBxPjF6WtzKysQ41g4nIlHQpZZq7e2c7l2xw75fGPD/ZMjo4pM8K/98aejfkuSpM2d/PlrsytrW4Op+C2HJkYy6fGYachYVOJ2CVLARCMjxjBGkjdFAGO9SgwvXGacu9SljBGCvZnk4SIKARTFBuId13UppYRIEiE33qQUQkBwt/E24I7jUJcSSSKS1IPvrutCCAghvRjddanj2oTIkiTBPcMEloDdbhLCyQjz6BFTjDFGqSTfGMY5d2wbQijJyt5IjLqOJMl7sjjAcRzAgfgKkR88vVo5+9rZ4yfuUBUFQsQ5oIzNz13O5XaO3HSzaZre90KwtZ31+4OWpQtai3FWrVVXN9aCwVAikezSuAgiuLGx2ZfuE5y3S12M0OLcdNtuDY9MQiHZhNCyrPn5mWQyJSsqgBByrppWfnt1Y20l3jcgaoQgQqYvUNzdrpYL0XhaUAmKqhuGeeW1Uy51AuGY6zgIIcMf0jTj/OlnU5lRiUgQAlXRkv3Dc1fOLy3NxZOZTsdmjGmGFU+lp86foYwGgmGCoKpqg8P7irv5s+dOcoh102y3OrKiZDL9pWL+2vSlQChGJCJLUqpvQFf1F597stRu+Xz+ZqUEiNTfN4AwunT5vG07fp9fkaRkMpVO9V25+NrU7Jxu+hRCSsV8PBEPmNb1lZXtnR1VUw1N7U+lx0ZGa9X6iy8+v1urqarerFcbjUY8HHOpO7+4XKiUTUOz/L6hTF/I8l+cunrm8mVJMWRV3dlcVTVVUpSNnWw2V3SpG/L74T+9vDK/unn+6nRfMnnTvtGgZTDOy/V6vlz7yG0j+5IBgWQQQoxx13U54ISQXhaJciZyFLDbFhtCSBkVKiCEPWEl45xSKkwIdNUiNyyBEBHccA4YpRxwjD3SiVEKIGSMcc48gxG0KWcibSd2y/aglYiUEPTEtuIKqQs4wEQSs5lRKuJpiLDQXHmomzHqOpKkdHUcnFHKGAUA4q4FiqlPqQsBxIT0gixKHcYYxkSgNXGJf/jvz798+tVbbn8AIeQ6DmW01Wy8duqpjkPveuC9iiwjiBDGAILrS4vJaCIQ8FNKKWMYwI3N1UvXLkWtwO133MsABxwiiKr18tLK2sTYOCaEMo4RIjK5/Norm5srowMj4wdvFaE8hGBpab5RLew7eAsAAIq9ehB4+akf0Ebl6B3vDMb6xL00K+VLp58YO35vIBCjnCMEJUlqNWuvPP19E7pH7n6fPxzljGGAVq9PbWfXRg/dqmo+BBGWiaKqtXLpwsuPE6dx4qFftMwAp8x2nbmps5TxgbHDRJIlWZYUVVallaXF+bPP+vxMYm/sAAAgAElEQVT+m+95WFM016GF4u7K0gyW9b6hfZKsaooqqwomeHFpYfbln6QGho6cuMfQTbtjLy3P7+7uhBP98XiaqIqopuSML81enTnzzMiBIxOHjvtVo1KtrG6s7W5vJYbGwtG4qiqIEEVWG83G7NmXl+YvDo9MTBw+Fg8nKsX81vZWrt5KZoYDwYCmqEQmEsa1Wu3iyafz+Z3MwNCBySNBf7BQLCwtL+P7P/bHmqan031WwJ+rNC5Oz167Nm07rmUYx4fjPhW7jturrcMCPgEoOBmxKTBGCEJAXddxHM45whiJyQchAIAy5oophUW+ErjUdV0bQIi7NXUi3qWUMuqKY4WXcB2bui5CmBDitSaCEABIKeWcS0QSJAjn3HVsxiiRJOGvPLKLA+q6CCNMiMhWcc4du8M4l2RFtI3qnhNQ15VkuceZcc5dpwMAkBVVhKS99wFnXV8h8lOMujaAUFYUQQmIwT88eVELxPszA6bP8vv9ls9fKm4vzlyxfMHb7ro/FAz5/H7LMjVdL+aLAwOZcCgcCPj9fr/l87Ua1aWlecLYidvvCgZDvoBlWUYgENzN5/v7+8ORiOX3Gz5L03VG2dryXKeSO3bng/5QyB/wmZY/nkwvzk1PHD5uBQKKrvkCAc2wNE1fvT5dL2wcuf2BaCTkD/hCsWg82b84c3H08M2BQMC0LN3QTX/YsvzLc1d2V6cnT9wTj8eDAX9qaNTQjbX5q0MHjvqCAcO0ZEW1fIFwvG/h6vnVa+f6Jw4k+/rDoeDo+AGJkFxuu2943LJ8qqoRIoUjsUjf6MrM5cVrZ/pHJjID/elkYt/4JGBupd5M9fUZpqFIMiEkEo4khg+sLc5eOfW0GQmNjY6NjYzs3zfRbtaL9VowEjF0VZRiRuKJvvFDW2vLl049J6ny6L7xA2Oj+8ZG6+VSoVy0AkG/6SMEq4qSHh7rHz+S3d4498JT2ztrmcGhY0eOHBofljCvt9pYIqauEow0TRsY3T80NlmpVC+cfnF1fSmdSt52/Ah+6Nf/GCJEXadSKmJqH9s3eNtNh6PhwOr6ylBQSQQtSZKIwD89AotzsYsKRhhC4LqubdsAAEmWsdcdBnR9AkcQypJoowoopY7dAQBIstrVOHgTlDGKEJQlSSz/LnWdTgciJCkq6tbdelOZUoyQYF0BgJS6jt2GEMqKesM2oGCxXEwwxkTQQZQxp9MCEIlopJeshgBQ6hIi9agzzrljtzmA3khww5Bc19kzEnLOXbsDAMCS4Ha6BCcAX/7p8yP7j+qaJr6LcTZ98Wyp4/RlxkZHxzxKEEGE4EZ2J51OKrLk9UBhrNZqrWxsyoo2MTFJiFhrIMKoUm9ACC2fT/wQEEJF069fu+w4TiyVDgUjCACMAMa42WzWG7VwOAaRl8G2/KHd7fX89gpW1ER6EGOIIdIsn2N3crvb4WhSlPUBwK1wFEvq1tJsdmU+M3ZIlhSEgD8UlhX1yoXTsb4hjLCg8lXdSI4c2FpdnDnzrBlJBkNRhGA4FPZZ1uVLZ3UroCiKeCK6bgxMHG522Mknv+NwFkukVUWNxePhgDF77SrARNcNBBGCSNW0gfGD/ljmwqnnr105ZwXDsUgsnYwnw+HlpcVCuWoYpljdVFVLD45lxg+uLs6ffOEpmzrJRHJsqD8TT6yvLa9srBNZ1jSNIKRpemZofPzorS4Hr77y3GsXzhBZGxvoH0tGEaQ7uXzLdiWJyIQoipJIZyYOHw9GktPTV18+9Qo+/v6PbW1tGZgfHekfTMVKldLzp1499dp53Qy+/eYDUZ/u5R661diQ8/zW2vNP/vSRb379a1/72uNPPYf9yYmRDCFSb5XNba89/9Tjj3z9a4988xtPPvO8q4RHB5K23eGcS5KMieQF3hAAwKnTefXkyURmUCFYoJ3i7ubpl579wfe++61vPvKjx366VrSP3zQpwB5n7Ea4AoDj2K7dmbl8XgokTV3pze/c1sq3v/rfv/jNn9z30EMKhoBzSt31pdkXnv7Zd7/97UceeeTpZ1+U/KmRTEJEKRhhAZAEanId2+00z52/nO4fFH5PfB9lFEKIMenR04y6jLoAIkmSbxgHAJzz75+azQyOCRGHbXcqlcrUhVMdgAcyA5FoVORMxOPa2t1JxRMQIQYg46DT6ezkslvZLCFSNBTSFA2LJAyELmXlWtnr1sM5pdS2O9mNtQ7gdrUYjmcwFuQHsHyBq5fO9o+MY4RFwtSxHULkbKm0u3A5FO9DAGFEMMHhWHxlbhqpqm76BDSFHFi+YKXplHLr2fUF3fQDjglGoUhMJmRm6rVIMuM9LggIJoFYOlcorlw5BYjsOg6ERDPMTF9mduqCA4Fu+LwsJYKBSBwbweWZq2tLs1YguLG2aliBof5MvVLa2t42fRaRCIIAIej3BZID+0ql8sLC3FZ2S5Hk1aWFTKY/YpnLa8vNtq3rBoQAISjLSjTZ7wslL1++tJYvtWynVS1Xy6WhTH85t7uxucExVFUNISgRHImlBkf2t10wNTOXrXVqnfbu2mq1XAj7/dVKpVxvcA5kSUII6oaRyQyH433wN//7T6uV6r0njlXazqW5hdmZqaNHbh4bGyGy9L790YGACrq8LXfaTz/23S996cuvnLlgRvtvPn40ErQun36Wpe556SdfQgBw2nnuJ9//8pe+9MIrZ+VA4sSJ47GQf+bCyzk09uqL31MgwAiefPL733/8pV/4+B/dfWycc8ao/a//5Q8+/Y+PPX/x2oG0ce38K1/64r/+5MnnGq504tZbBzOp4sbsY89dv55biUkAIrh05dUvf+07I7c+/Kv/ywNCJnHysS999Lf+9FNffPZ3f/EO5nZOPvv4N/79Kz97+kVOFKYnz09dCKPWk49++ytf+eqpsxet2MDNNx+NBKyLp54Gffe99OP/wagLAXv20Ucef+HCh3/7z27e30ddh7nt//s///bfPXLutWuXhyIm7ApCXNeWJLnLV3POmWt3AEQCdPXWdQghpfTPv3MGq/56rd7pdDBCxfLO6RceR2b07Q++W8bEtm1JkhRdQwRPzc4fntjnOHar2XJsR1WVWqP+8plTCka333zCbwVs28WEqJrScDrLKysT+yZbjWa71eaM6ZZZLRdefukJXt5+5wd/yzD9tt2RCEGSdPHCyUR6wBeIOQ51Ox2iyIZl1WuVF370VVjP3/OBj8fj/W7H4QR2Oq3XTj9/6Nb7OCS047iOK2maZpqddvPkD//NruZuf89H+vsnHLsjEWltZWFzd2N4/zHAYLPdBgDpfp+mGbXizqWnv22Xd48/9IvjEzdR22WAT10+T3xWMJSglLc7bVnTTF9AUdVGpTR98vHC0tWjdz10+PidrUbTpfzKtcvJdAYrBmOAMqCbpmYamMjNZm3u/MsrF19MDk+O3XRnIhwrlUuLK4vhcIjofswhJLLh82u6LhHSsTvL187Pn33OH43vP35n0Aru5HI7uayla3o4BQEyDJ9umrIsE4xt116bm5q58BKEfPLILdHkYL6QLxRzEoe+eD+RFdOyyNM//m40NRDpy8Qi8YMHDoyMjpdr9bmldcbYvWnVNTEXqgkIf/joY7/3+5981wc/9K2//PwdNx+UJald2Xzo1h+9873vLmXXn3zse1/4p3+a36w89IFf+uqjf3PHzQcJBNypvu+um9/+y++n9eKjP/7BV77ypTNXV7FdMUbuvO3QILWbn/+LP/zcFx7JHH1nJsD+8nc+9K/fe/7Y3Q9+7p+/+fDb7zV1BTD3//jN9x978GGtVXrxmee+9c1//8ETr2gSHFu1P/Lee4hEnnzkH3/j9z/VUVP333ngR1/8+8/+/ed3avSh93zwq48+d/XHn//+nDL7/Hc+/anPLG433v2Lv/yd//qFW2/aL0ukU9l64MQPH37vu3MbS0/++Idf+/q/Ty3u0GY5ffxdR8fidqP43z7xO//8yM8Ovf2jSRN8/r9++v6P/tGh/gh1bYgJFx2vIQAAOqIGDULhEEBXl0UpdV3HaXcoaEciIUwkl7G1lSlEFALccCSiqSoA3HVps9naXLqe21zeNrRkX8YX9xFCOOAwX4B2i0kSISSeSHAIHUrbjUZja3Nt/mosGg2H44FQSCBA3bJkzh1VX1+ZufOB9xCEOOX1RjUWSV58/sd3ve/XAuGQ6NDDIVA1bWDyxNKZn114+Sfv/difhaJRCHizUR8aHn/1J9868e5f8cdiBBMEAIdQUbXj7/jIq4998cyT31V/4eP79h2RELT8Frjozpx66vDbPpiIxrtomcvJvlvf/xvnf/LvZ5/8/xqV4h0Pvs+vafFY+PKFs3MXTx2+9x0xrQ+LbZ0glMPRWx7+5esXX7l48mfL81fe/gu/um9kKJWKn3r5ud1S4eAdbzdNfxcDI8vyH7nn4b59R6aef+zkY18+fOeDt9x+/+BQ5pXnny6vrxy4+e5gKCLksAAATVUmb7pzcOLo0vRrZ578kWLpt93/8PjYHU8+/mO2vT55/K5QJNALfRVZGjl0rH/iyM7W6rXTz02ffWn/8dv37Rufmppq7W4MDI/7fBb80+9dsHyWTLDQLlHGOQDtRmtpcf637t1/YmKQEEIppa67lc0h1RxIhrq6NfDov3z6I3/2/9xy4uj89FSkf9/bHnr4d37vd4ZTUdexAQCEyCe///l3/dpnjt18fGXuqi8x/OCDD9x608Cf/tnf/uTV14b1xid+99dfnCk6u0sP/dqfdq6/cHKx+a9f+uoDdxxGXbBUXDx14Mi9qYmjrfxaC1lve/tDt91+7F/+yyd/+x++/7G3H/rnz/2n/+tLj8cDKLj/gbeNS//89Z/+7p//xcc/8qG+eBiwxjuPjZ9fbUia7wMf/tgn/uwPBlPRHgL60Rc+85FPfP7EiSPz01ejAxMPPnDfodHIp/76fzxz+pRRW/qPf/i7U1laWb76v37iv22c/N6Vovq9Hz06nvAx15EUtQfkGGNOp8UBlCQZCyV8F2AxxlzX+eLZXKlDRZ7ddp2ffvvf8pVq2B9+74d+HWOMIOCQcw6r1fKLL7780NsfUhSlS7+BQin/g+9+A8vyXbfdvf/AYe/EgNuO+71Hv3ff3fcFg1He3TaIMnbmuZ8sLc8pbvPDv/MZRZYwQoxz23Ge+O7Xho6cyAxNiJ4jAic3G/XnfvDVxsbUxF3vu+tt75eJhBBwHfrKUz9wiTJ54j60p+rY5WBzfuq1H3+ZSOS+D/3u2NhBCSMGwOzFM0vrq/tvf5sqeZEG4IBy3mnULz317e3ZM8n9J97xwY9FQmEI4fri9VOnT07edp8/EPbiN4FRGS9tr55/4puN0u7xB9533wPvMDRj8frCyTOnosPjfUPjEsYAYOApZbjrOmszl6df/okk4Xvf9YuT+4+sbGzPL8y5CA+N7jMtv5BOAgBEZ5ZGs3n9yqvL0+dSmcHDJ+7eLZSa1WKuWByeOJxK9WMsiWtBHHIIHMrKhZ35i68Wsut9AyNKOJFM9ZUrNfze3/6PAEJKmcsAY7xer09PXVxanNNN666DIzGf5roOhJDISigUCFp6NyoBAIBWrbhb7tx6z4Of+eu//dR/+sS7Hrrf0mTmuphIkqwgjO1WdStXv/Xut33ys3/zF5/+5LsffseP/+1vO/FbxpSdj//ax5vBQ1//8t8/9s2vvfrqqejkfd/81jduPjDUm4IccKfdXFrdOnD0tt/7xF/89V999gPveWdh6qkfXqh99J1H/ug3f+XZq4Wvfu/R0vQTTz39/GZT/9evfeujH3go6LMABO3cwt/909c/+PE/+cK//L8f/uB7Qn6z95MDAJu1Yq5i33r3g3/5ub//1Cc/8a53PvTNf/jP1uRDVvnqb/1vv6ePP/Ctr/zN1//liydPvTJw4l3f/MZXhmM+17G7UbsXqzh2hzMOMSayDG/UEAqGgCJEXtusdVwuZnCt3jj/8hNED6TTAwMj4zfCMM6b7Xah1hjqz4h6RogQB8Bud5aXFolmBnxmKtmHoVefjTAu1tqIueFIbM8dAcb50vKCXdwMpocCgRDBBEFEENKC8SuvvTwwuh/e0KQBLMmSom0uzZY2rscHJzVdF6xgPDM8fe5lYvosf7ArxIYAQisUBUTdXbiysTgTHRxTVF0iOJbKQMeeuXIu2jeEMRb1EBgCJEnRkUmHgo2Zc0vXrwZSA7pm+H3+RCJ1/tQLnGDLH4IQiGoAjKBq+tOTJziAU2deuL4wE06k+vsHDCvUrJfnrl0xAiFN1SBEQiBLMAnEEoMHb3U5P/3cTxdXlsbHhgf7R2zX3VpdzBfylj8gYwl2hV6KrMT7hgYnj9cbjdPPPV6qV4fGDozvm7x85sXZ6XOKYRqmX2SjEYCEIMOwMsP7+8YOV+vVaxdP1xrNVF8G/tVTiy5nlNJSqTA7dbZebx49cQej/OLl85/9pfvvOjIpAuteeqGHJcRKKSgsSqkQm4jGaLCnD+0eIeSDnPM//IVbv/HMtUhy8Df/6M//4Dc+pMlyIbteZ8pQJnVD+s45Y5RRJkoaxAwQmbtv/J9//Cef+4ruC/+HX//9v/jkn0T9Wr2cW9upDA30yYRIksQ4Ext+tVtNIsmCKfZUbzdEX8yxO7KsiMw6pe5H7ht/4uJOrG/kjz/1V7/xy++TCc6uLtrEzKTiCALXdQCAkuiKK0QujFLXAQCKJHpXgthNbtq2LMv/eHKj2HTqtVo+tzt/5ezS7EUplBroGx4emwhFY6ZlCSVSvlCYWVi588QxjAnjvFatFvO53Z2tuYU5ohlyp3ritgcCgYAvFCBEBgDMrW4WdzaO3HQz4Jxy1qjVCrld1+6cPfOcXcn6DfPg8bfFEulgJKIZJufsx499Z2T8UGpgBEDEOGs36vmdHcdxdjaW1y48YYXjmeHD4/uPmoGg6feVS8Wnf/StW979S4bm1QZ2Oq3izk6z1YRu6+rz3yO6lukbGz9yZzgcsUKBtYW5K7PTN93xdkVWEUIMgHanWcxma7WKZvkXzj5Vz60PjR/GkjE0cTAcCl25esWGYOLwbbL4UQC0bbtUyBVyOdU0O9X84sUXopGE3bFTo0diyfji4rwSCI1NHCKSggACAFDHLuby+VxOMS1NIYuXTyG31SjuaqFkon+0XKuGk5nBwVFZkhHEAALqOuViYXNzGypyKBov7awVN1byS1MtpwUUIxhLTBy5Pd0/rMgaBAAi6LpurVBc2dxgiMRSacQZ/MzjMzvbm7NT55YW5xqlQjAYG7v57nAsFfCHP3Zr3/5koFdr5FkHB8I2OPfoLZEAQZiIuS2ISW/GCJEVo0JTyRmr5DaWN3Ij+/YHfKZI/AEukL0nHBSMqkg/cACo63BRjC7JCCG7VZuZvR7rG0pGgz1v47qOUK0L8aAglBEiWJZhF1p4IlmPye0I6kkIQp1Op5Bd29itjE8esnQVCPUi9CrNOGOu48iKLITaIh/qdNoAQoSIJMviLjjnCCKAIGeMUipJ0mcfvbSWK/l9Plkzv/vFv+pQhMzo/Q++J5lONcqVeqWi6Jo/ENwtlda3dk4cOVAuVdqNhuX3+wP+5aWl1869wlWdFrc/9LH/HTNeLpZs1/EFA4V6c3Z2+tZbbq+VS/Vy1fD5fKEgQPjVZx9fX5unuwv773z47gfe1yiX27WaYlrZUm76wqk7HvoPrVqlWi5pummGIoiQVrPx0g/+rZVbVTT9Ax//c5/pL+cLCOOt7ZXlxdmb7n+/3WxWiwWsqL5QVFJkTvn6wpWpZx4BrjN69M77H/4wbbZ2dnfKlfzS6sJNd72L2nYhn6eE+MNRTTMgAK7bnjv5xObUKwCCgaP3Hjp6t91uV0u7K2uLk7fejxGpFooOZVYkbJo+hCAHsFkuXHnxsfzC5WBq4MAdDxlGYHt9ZXt3c//Nd2mKVimWHcp94YhlWV6TVUZ3N5ZmXnmiuH09EE2lJ050Ou1qtTJ+5LjPDNXr9WarbYVj/kBAwpJY4jud9sbi1PUzzzQKW2owjHW/avhHDhzzB6KtVqfaaFjBcCgUkYkkmvTilj8xdeFkdmHaqVb6Rg8dv+fhkdHJWDhkqMrRvmDIkDn3RCWCbXUcx+sIzyjnHBOJSLJQkUAvW4YYYyILLrRPAECEEKMuo46iW+m+jK6p3v4G3VbQTGghOXMdG3ncK6euLer1BGaDEBJJiSdTlq4y7uW8qesgiCASO9Nzx7EB4BBLXfDTq4KETKhKXKcr1kIQQddxGXU1w5dKp1VF8QxDCAY4Z1SMxz0RP4DQsTvCpRIiQQGNusE788SRCEF4frNhBEKqqtZqtYunnpJ1P2LOoRN36ZqhG7oVDHCId7Lbs1cvOpRLAARDoVg8rpsGRLhaq26ur1DOaLsycfC4ZZo+v183tXajubG6upXdAK4bDkcjyYRmWlBseeHaG8szwHWcZmPi6O2Wz+cPByHgzUpleWWx06gGo+lwPGn6fMLJY0kisrqzOs/cVrlSGjl4cygU1g2ddtyFuSvba4vBxEAknrL8AVmShXbOCkURVopbi8WdjXK9se/IcUaB6g+WsptXXnlCTY2GE+lAKKTJitCmYUzCfaMAyaXNxUp2ueM4mYnDwXCsU6ucffq7FJHk8EQoGtN1nWAsWl9LqpYYmZSMwNb8ha2Fq4rlHzp4XCHk3DM/2Flf6Zs8Fo+nDE3FohE3gghh0xdKjR3WA/HNpWvF5WlZUZLD+5amL1w9/UxocKJ/eMwyTElkphFCCBKJ+COJvv3HjUhffmOptb2CMcqV8jOvPotVfXD/0XAgoEqS6OmKIMSOrHYqxdGjd93zvl89cPz2WDhiKIRgBACYTJhB3UseC2TCOEcYc+pyRjGRJFnFWELdjay7ZKdXDuE6NmNMkhWR9OCMYSIRWe2q/W4UaHgMqetS6sqygjCm1HXtDuAcYSLJCkS92g8Au18CAKeOLQJlBCF1XdfuAMARlqSuPsojFTzMDqljI0wkSYYIAQgdx6WuDQBAmGCRzwGvO0TsIiXL3ngOAHVdRh0u9ruQ5B646uJ22M3NowvbrZbDXEpXV66vXD2N9KAqyQeP30EIQhAjACWJmD5/vpCHRDp69CZVVRCCIvFfrZaWFuc6rbZTL40fOCoKCRHGqmYEQsHp6av7JyaC4SiASCicOedElpcunwEI2+VsID0SicQwRpKqhMJRl4Gdlenhg7dKBHcfCwAc+AKR/O5uM7/ezGWZrKb6hyVZCoTCyf7x6ZNPhPtHLX8E427FNYIQokAiQ227tLFY2lzIl0uDB45qupUeHNtZvV7YWkyOTcpERd3yZIQAxiiYGtB94d3la8WVa7nNlcjA+PD4pGqGVqde5ZiEYymCRWW36MYACZGCib74wER+fXHltecK26uZA8cjfaPF7NrGzDl/NGlYfoi8rvdCSCpJciiWzkwcb7U761dO5ldmo8P7ffHB3MpMMZ8NRuKKoop6LQgghgghLBESiCQGDt0qmeHCyrzTbmmxVK1S2Fq4yjkzraCsSKIxAD7w8K/c8e6P7D9yS8hn6TIhGDDIHcZdCg4krJBGGGeuY1PqQowA50IYQmQVe/oOsOfFPXaFuq7rIEwgQow61BHiP7WbK9xzkIBujLtuB0JIJAlC5Dod5jgAQizJEpH3ztvu1wDGXOo6mAgeCbiuQwW4IhIW5tENTHsvYQySLCouOKXUtTucc4gQkdU3HsI5B9x1nK59esSRY7c54AAgQiT0pkaMoj5EiMrOrteatmtTfvX8y6X8th6IR+KZ4fH9ossT8FAr2NrcCISjqXi0J0XgAFRq1Vw2y4gM3M7A8HjAH+puRwUxITulKsYwFI4B0K3ig4DISm5jtQWgUyszzscOHO0KYIDPH7hw4XwsldYMy7MOT76D9GB4/fo11qkUN1eSY0d8lo8gpOt6qWXPnX8hNX5IluSu9sBbowLJoXq50MiulrZXKm071jeiKLJmhlvN6trc5cTgPkwwALyLECCC0IwkffGB/Or1Sm49t7YUTA0l+wZ9sf7i+sLG2nw4NUAkqVdmhhDECCmGFR+7iSOytTC1MX9FM63Bw7eFY+nLr/ysWq+GImlEcE/m4bWUl+TowL7Y+NFWs7k1d4k6ncHJY5Y/MHPpTL3d9gdDooQO7qn/I5iE4n0DR27XrWB+bcFxHD0QrVeLq/OXW52OYQYwlvBHP/svkYBfVwjBkHHgMOBQQBmnjB6IG5YMqeuKMjfOGIJIklUsSV3M8Ubr4Ix1qV6JM0apyxnHskwkBXXlKF3T8MqZKKWuaxMiQaE3cTqcMYiwpKgYE9AVRPWqwkW5LKWuqCVCCLmOTV0HQIgIIZKyZ67z3rVR1+EAYCJhYeccOHYbcA4glGQFQdzzBl1bANRxAESSRLyqSc4pdbnrAgghRJhIr2ewPJUk6u5td3q9WihV1teX5y68bEMZEDUUilqmqZtWd59aCDhYXl0NByORcECIIznjpWJhcW661Ww5AGFq03bT0EzNspAI1QAvNzuNaimR7OteMWecV/K53a31eqPJaadZyspGEDGkmyaGSJakesfZWLyWHhjvyREAhK7jVHazHZc1ClnmdPKFvEs5te1QKAyxXKnXdldnkoMT4ofjAhwgSB3HpgCqer28U9tZb7n29sZms1YePHBzs5Jbmr2QGBwnRPb6V0CIMEYQSqpBsS75Y8Wt65tL1xTdquRzViSuStLVsy9EUoOKqol6Qy5STAgSSfZFUm0gGdH02tSrjcJGNDWs6L7l2Qtr1y/5ownN8PXWWwghRohgpJuWpPmZGYsNTqxcPduslJL9Izsrc3Nzl4mk+vyhHm5BgAuFjiJLgUgiEMtU6q3k4P5Op80BqtfKs2eeKTWq+F0f/xOCEQPAcZlLuUOZw9xSuXjq5LM3pXwDCS+NgBGBEEmS3CXL38I6XMcR1DBC2HVtzgGRJIh6FSV7PYdXfei6DqMUQiSCFhbN6UYAACAASURBVOo4EAAiK9DTOO3loERcLmJ3SiSZMcoZZZQy6gIAiKSI7mYCNO+5NkApZYwSsdUdY67rUNcV5iEsqidP7k45IEIWWVIggowyzhh1HeY6ouBV+DrOGLwBMD2/JBFJcAA/ePFytdq4fPaZ3OqsHh1AjBm6Fc8M7KytYEJkVRXPbX1zMxaLB3wWALzZbK4uXCcIFvPZVrvpACwBVlifP3jLPYWNDQCBrKoQgZbtZLPbfZl+DgFjvFarblxfkBQtEk0szlwkmuHWC4X1hYljd1d2dingiqb4fYFzZ0+mB4ZkRRdFbqXs9s76aijVnxkeX19dZJ1Gu5bbWZy2UqOVUsVQpGBiYOnaBcpZMJYSyxR1nZ311Z3sVnRgLD56yG53qvn18tZKaXlaDUYwkSPxfrtVW776WmxgDBMijnJde3v5ejabTY0c6Bs9aIYS2YXpzYUrucXLzXrVF81EwvErZ54nuunzh7xYD3Cn01lfmCsWikOTR5ODE7Ghyc2lueVLL+cXLiqygoi0OHOh1WwEIkniLVWAQ1CrVuenp7hqDIzu94ejqbHDruPOX3ipvn7NKea2tlezxYKsqIZhAq97C4QA1GvVuekrNZsNTR4LRqLJzLBhhRqlfC27Urx+ET/wK3/oMmBT7jLuMFapVi9fOXf2mR/vzp5//713DPalb9QYYcw489p7dedFV/7tuo7DGAOccU45Z5hIwm+IIifGqDiGwxtTUHgbCCGjLmdUdECUZBVijCACgIvGInuryV2nAwBHhADAmety6oqKaCKryNOoQ8bFxkBdOT2jjDpEkgWfxihlXqM3gIiEPSW/ENjzrlfgrmNjIiGEqEsRQhxw6tieKSAsIhlhJIxzwXp5Unns9SCcKtA2kV576WcOtY1YBnC+7/CJvr5BXyhcr5RzmxuypiOMl1dXE7G4okibK6utZjPV328FQrlisdmsd1xXleVGrXj0tvtD0Zjdau1ubUmSxDFZXFpM9/U5jr2xeN2lNNU/pFt+xbKW56eBJINmzaVupH9seGLSaXdyG5uGoTdcvru5HE8P1ivltaUFzfTFM4OyIhNJRpK8s34dUJdy2mk19t96TzabrxV300NjV888G4inVcNfyu9sri4boWisr1+WCYQwlBmtFnOtcp5jVC1sBtNDgWgKQtKuFVfmLkcHxxDC+Y219ZVlK5pK9g0omoIQ9IXjgURmd33BpU67VnQalcjIAZ9mzrz2Qtt1wrG04zq766vrq2vBeDqe7lNkGSGgaHpy5BDHUjmftZuVTnGTSErH6SzPXpIMn+UPOY69NDezWyqnBsbCwZBMMIZIIpIvmkyNHmREbdYrvLLb2FzaLedz5ZKm6bKqtRrNpfnZbL4Q7x+Jx+Oa7AlvZV2PZoZD/fuQ7seDd71P1jQOYa1em5mduvDKUyunnyROJzZy6Bfe8bZMPAK9yAtCCISjp4wJBhZ0YRVjjDMKOIMigpUUhEg3fBAvxBhjnAk7cV3HdWxBWHFKxThMZCLJ3i7m3jd6tJiYmo7dAYATIkGIqGOL7sgAItLV6kIvir9hXRww17ExJhBChLFwBSLm9kJtYUpQcMGQMQoES+Y1LIWC9HJsuxtkQYKJh2hFqCisizGxe5twYgijM+vV5fW1ufMvAUkmkqYQeXTyJtM0CcGGaamWld/aXFteLDaawHXtRj2RSkfiMRHD7O5uV8vFer2ia2qttDN55BZd0w3T8AX8xXxubWmhUC1Xd3e4SxOZoWAkQrBIPPNmtVrYWmYQANphAI9PHjV0wwz6r01daTYaSwtT7Y5DiJTsHzb9Ptzd79wKhHc2VjuNEoSgVSuqZkAPRsPJTKfZrJRLi1dPN5s20az4wIhpGBL2ngtEONI3mt9Y7LSqnLHS5qoVTyWHJ3XDv3X96urM+Vq1IVuR1OCwaRgEi/JMBCDXfOFw/1hhc5XajVajWtpZS+w/Foqlr597aX1pOpvNGaFkemBIN3QJE4yg4K0QlkLJwWBqqJzfYYyDTt2p5KVAeHPx6ubCbDZfiPWNJFN9qiITImJkT5WNJSWWHgn3jdRt12nW3exis5DdrZZXr11aXV8LD+xLpwcMTZEIJpgQJOhJBCHQDCucGsTJ+37p7Knns5ur1y6fvn7yidb2SmRg8uDd7z1y54N3TvRFDMWbd6C3Lnt5X9dxqOsw5gLOOKMQQogxlhRMJNitTd1DJwExBanrUKfDOcCEcEoBYxAAKBTpXkWhRwoBz04QRJC6ruvYCCHBjLm2LXgGL4oQlGvX3fQsjDFK7Q4mHk/Vi5GE3Uqy4vXW20ORiaSN69qEyEJthRFyqMtcpzeGeLG+90TERXLAGXUxFr8MAgC8ulq6cOFMdmkKEpm7/5OvN+uOLEnOxMzc/a6xRyAQAAI7kHtWVlVXdXWzNzaXZk9zZkjOAw/VR8ORRs8a6kGPetbLHOkH6IXUHOkcSuKZEcUhh9Ncem9WV1VXVVZW7gkkdgQigNi3u7i76cHvDSCri4ODk1WZwPV7L+DmZvbZZ58p2/XvvP624zicAUMQQmTyJcuxHz9/emNjY/P6Ndf1Ev9KdNo4bZwcjIddRiCH3ev33slmspwzLoSfzTm+9+Thg2p17vrtNxwnBRsBNCGR3Pv058z2MA7G/U59+14um7Ut4WUL2VL1ePdZxrU2br/t2Ea0iiU9ncjyxcrxi4dMRqjk+dGuW16aW1jJ5ktz9dWDpw9oOth441dcyzKdO5gObuGWValvtvaf6nAEUXC+/9SfW5hb3lrcuLH/6fvTbmPt7juZTO5K1g6ccYbketn61u3e2WnQbcbDfuP5x15lYfvNr7346Meq31y+ca+QL4m0XzW5liECutni0vXXdRz1GgdyMgxbR9nKIviZwd7D8uJyoTJvW8LgEyy9ykCttpdb2Lztl2u987OweRgFE8qX42mfk5qbX3Bdj18elQbvYgyAAPjy175zcX4y7p7395+Qkne++Xtf/Na/qC6teI71Zr1Y8q1XE45UAE5JrSVjzJgHAHJhm7N85nBmodHsWq2VlhEgMsa0jIEUADAuhO0gT3PlK6X45Lr04LdsW2stoxBIA0La6cFfecLZXYlkHCFjwjJjh0jG6YWAl24HPnu1Siro9ozKbnyXqTFzYZljPiFlzMr0SgGCJSzzAwCifzjo/eBv/uN00HWLNa3U/PL29o07Qsx67gkQYqmOj49vXLuey2Vn2IcGap41OudnsdYZz58OOxs37hWKpXTiB9mOO4iUHA+W1jZeUZMAcB1v7+kn3HbicEJRIIW9uX1TcOa4VqR0exo2nn+ycfvNK746Qam8bGE8HHUuTgkIwqmKpovbd5iwHNsJFbR2HtiuX6ktG8kAxjAZ64tkOZlCtX768pmOJioYtQ+eFZbWS5UFhfZk0G7uPKht37FmDWeXVTAQllvdvB1MpqPzYxWM+kc7JMTc9ptRMD74+MfuXLVQqs6E1mawmKmBlJa38wvrveaJjMYyCt1c0astHT7+xajXqSzUhXBMZ5vhqpjNzhgCQiZfWbz5Bae0MB70ZDCOCYeT4UXzWCtZKFYYF3Qpbmh4MYyruTpEoQNs4+7bX/qn313Zvu25rmsJV4i7i9mSb832nNkLWisZR6Yv16TXyLhlu0xYsyjnqkWlJBWScaSVZFwgMq2kUQHjli0sOznLZhv2EoICrWWSEnAOyS43wQ6zHAfxl0Y2p1fLOEJEnoLFpgnRJELJLr+EvC4vNIQSJixjP4yhlJKkpMSnJUT3z4OSZQJJJLpV+P0njR///V9IZPnqmoqjtWt3FpdXTCkNkqMGRqPBRae/sbLqet4Mk9AaWs3GeDSMCcvl+f6wvbS2NTdXEwmYhYQwCuJm43h98/oMAkEAAo3C6pyfjUYDqTVFQTjsXf/CVx0hNME0kr1BfzgaCQal+UWWQkCzcylbruzvPJHBkCk56Z67+WK5tkakwzCurKw/efdvaxs3/Ewu3ejJ+cIYc3MFxy+evbgPWkspu43DysoGab6weavd2DvdfbSwcetKVyYgAmcIyLiwqivbCnnn7BgQBu1T2xI3vvSblpd79v73paZKbZmnuv7mTVNxVOYX5xZvvBEr3e+1p93zaBoUl69Nw8mL++95uWImVzINauYP06tmSoyWcEqLq8vbr8XRZNg6Q8BY686gf36yxx1XyYiZEh9RYiGla28srmy/843f2rj1mu/5Gcf2BLM5csTbC9mibyWlASDQl9ATAAFpADDtyPhLriPdc4lsgglvuBBGRAgAkHFhO8lOnVUZU0s0ZRKlpIpjxjkXFpFWsRH5RGDcunQ7gFewNWOOxoaNz0FEJSVpiQhk8iRhpcpxl4hwwh6NImHZkAJbWidLzQI+dlVSc/aaRi/YtA+DadhS//t//sHTT95nTsZysyglArqOWyiWkp5+ACLqdbvtdn9jdcVxHbNorNXBi2fPH32oFYVRJBibDDuT0SBv+9lSUTCBCBqo0+vv7e1c274huJWOHKI4jk93n0+DYatx4Ph5OR2oYDIJotFgvLBYU4Tddsctlg8e/nztxhuzJmQERILJeNTc280V5zrnJwSKCat7ceb5fuNgL4rD1a1b0yjaf/T+8rXXZrULls6lmI5H3XartvVau3mEgkVy2m4ckNbnZ8el+eXB4OLs5aOF9Ru25RIQIDBMzQshjsJ+r7/y+tejcBpNh9Peef/iLF8oKcLm/rP2eaOytGrb7mxjGesUHBljSqnRKFh78xtutthvvJz0zjy/4Dr2iw/+rhvr0ty8JSyGmHCOzH0RTaCotOr2+rVbby/WN8bdCwqnY63P958dfPD3x62GU6jk/Ky5Hb/2nX+1ffNutbZoc+ZawuKMATBERXSrlit5wqhXyShWMjLujkghorBsZIISvUP4jHGkLgeklFLGQJohGl6JCeW5sIEoVaiGhPdFl+5DyVhJidy0CEqjwAAABiXThgB2eZzPLgQlY6MdSppIK61iSjExxriwHYM1pXV6uHohIONCGH4N6dRlpQ7EhF6kNUuEs5LCn1YS0pzegMuI+G//1/+lPY0yc3XPdn3Pqy+v1xZXzvZ3M/mCsIQRpbxotQbTcH2lblkWIE2n08Onz+YWFo6ODy3XDeM4m83FcRR0mm9//VsXx8fCEpbrMIDTZrPZai3MVz0/Q4ia9Kjfa+3vVRYXX37y/ngysrNFGYxQyeHZwfzNL3Quuo7QwzAuV+YP919ms36xND/j2l2cnnSapyvX78zV6o2Tw3DURQAZx2fPP4rG/erKtcmwt7x9+2jveTju11Y20xIVaqD26Umzcbh647Xy4ppwMueHzxnpKBgPGnvT80OynMr8aq9z1jraXdi4yYWNNJuoQb1W82B3Z2H7VmV+aX7txqjfGffb4XjQOd4Jz4+4ZYcyPt59XKrVvUxutqPMbu+cHb3ceba4dbNcma/WN0oLaxenh8PzIyRwLNHdfXDc6bi5Yjab40lAyRiAgSW7zbPnTx/W1m/N1xYK5bmF9W1AHnQuGAMlo9Hew9PDF1NgXq7o2Db/9n//P580Tvuts/pC1RYCgRRgqHWg9N3FbMm3lZQyDkErZBwZEmnOLS5SRSlAM2roSjEheRUiLWWslQR9qSHNzPHPknDc7HuW0vpn1iXjWGuFDA0KnGruIxc2F5YRnzdKdFdV3ghAqdjIWyXXKnm5LjKTnSd6RUrNKidGmyvV+DFkEyOxpWYXc8552mls9BcxLTAqJZNZbURaKSGE1vp/+3/+vDeZutlyEIyzfmF58+bi6nqmWGjs7WitbD9LQCcnJ4NxsFZfFJbVPjvrNJpr16+7fubl/ksZREEc2MJSMpwE49e/8NXFer3TbA67ba9Q7PX6572eZ/FKdUErah3vB8Ph6vZ1z8tI4p12U2tCzpQMCSFbKM+tX9/deTHtdyvzCyTsw6cfr127yxhTpI9fPEWG9Y1rnAsUIpstHh6+AFQcOVpWFI6dXGFx7WbneH9p68azj37qF4qFQhUQJKnjZ09ipVa2blm2BQSlWp2Ad1uHjFkoBDGcXjQK1cV8ZeH8ePf89KC2tm0mAiolj54/7o3GGzfuZjwPEbllza/fIkXjzilwjrZD07GeDtzi/NGLh8K2C5Wq0awl0i+fP+wOxqvX7mQyvrE3P1OsX3tdKt093QPEUnVpvP/47OjFkFguX7Qs26TssVJ7zx61+721G6/ls1nBGWPAuV2uLlXqa2EQxGGUrcyPDp/3j19cDLoxMv5rf/hHlXIlkvr540fZfJ47TkwklQ6j6HbVK7vMwDhMWADAGBNWgh0ZwMg4TaWUESOFdGqRUkpKRSoGSsaggUnKLWeWW5pwlrQZaYBpTZDiOCTSaJqPrkRQiXmk9zYHebpZcUZFQca5EERaS3mFq4LCdoz6ThoQGvtMXJCMI8YFGrU7IRDRsFQoPbaS2CwpFTPS2kRflMw65Ea4CBnjjEkZ//Ff/PVA8lJtJZiMllY21zavZf2MbVv5yly/c9FunLq5wsnJ8SSM6ovzp3svLWGvbm9awtIE+0cHlhBhJD0/wxmMu+e3Xns7n8vlS+XTs8besyfM9gZBpKaDam3x8MWTXKZQW1vj3NJASsad5km/d+Fm8tF4gCTDYLK6ddvKlrLFUuPl81yhcHiwMzdXE5Z9+ORRuVafW1gUPGnH9/OFfrszuDgFUqg1EA3OTyur2/OrW/1GA21799P365t3tNYvH33iFysLK2u2EDw5LbFcq4+Go8H5MYE26Eb//LSyvJ0r106f3e+eny6uXQ+DYO/Jp06hXF/f9lLogiEi45XldeRut3FASqOwkPT04tQr1xqHO9PxqLywHEfB0wcfCT9fX930HFukHEbGGBNWdfVavlrvnOyPeu1cdUG2zzr7j84nY+FmPD/T73Uff/Kh5efXNq95jm2Z4kcSiJCwnLnF1fz84mg4cnNFNeyNT571+x3+G//1H9mceZmMnS0+ePhwPBr4ufx5r3P//nvvrJSWy3lANPMXhbC4sC53N87gX0CzUbRJUUApqbUiGQMiJnNiUVhO0tV1uUWT0AcAlDTlC5AySrSXZxMGERGRW3baeXIZXpkvme4UApJxBIiWZRuHMAuEAJLs/Ap0leQ+pLXWirTWWie/Jc4BQKnY0BbTZ2SX725embFZZm9GUyagMyIiyDj+43//HwdB7AgrGvXzhbmN6zdt2+YcBcdMvkjAH33488b5mQTsNA4ty79591Zi80S7uzvjzkUwHZKMUclRr33t5uuVclkw7PbHyvaPnj+ayrjXOtFhvLqxXapWBePIQBMIYTVOTgbNQ8t2ZTxBrWQwyc+vFOcWXd/PFkrt0/1pGDd2HyGz1q7dzhcLCTU7pYoVS5XjnadmdjbjDJH6F43FjTvl2tKo124evjg/3hkMg9Xrt+eq84JxU40xDEfivLqy3u+0g0mfc6NAif3W8dz69WJt7ez5J6eHOxfd/tr1e7X5RYtzxiAdBgOcIQIrL6zmK4uds0OGitmecOzJ6b5dKITTaWP/+enRYXXzTq26kHFtwWeTYAAZGppgvjRXv34vCoPBxamXL9G4Pz581un3+qPh7uP7q7e/sLSw5Nm2Ebzgs/3FEqzM9bJzyxt2phgRxMNe0NhjgqNAtAUr5DPbt1876fR/9JPvf/Tj75189MO43zZbhnFu2y5L5TleScjTI9lIRcVhYDArMqguMoAU7OJ8xoJN9+kVZ8K5lLGMQgAkrYx5mACIrniP2R0BZu4BGedaaxkFiMyyHCJScZSmNARm1J0QV5KOy7yPcW7MEhkz1QyjDz2ruxMAAhgW1lXTMlcjMqUUJtpwJo1kWhNpLRgXqMNgxHSEHBzHTis9yBkrlEtzq9ujTisctle3bq9vbfMZDxQRUQ5H7XAyGI0Hk2jCUF70mpqIIVSrlXw+v3brDTUdOK63tn0jVyzwRLgVENH1fNexQU1lPOWAAlHo+HzvoUYAANvxlrfvFBZX+51mJus7nssZE8mANMYZ48jylfnNu+8w0qhilBLjaHJ28Py9v4mV2rzzVv3Gm93TPS6HmWyeMWZaIzkyjsgZWow5jv/Wr/9evrBAcUDBVE9Hsn/+4u/+DBkuXP/CuHU0OXjAmEYgZKSJhqMRInLGOTLjE2obN7/wrd/nIhsPetGgp6Pp6PkDCMakZfvpu6rXSLXT0FwojCEyFIIDkO1lX//m79756j8Nh8N4OmEyCs72G0cvWcYbdE5JS85AMGQMGKJgLPlMzA0sxueX1m9/9Tv1t77FM2WmSEtESRDG8cXFiZqcs1FbT4ZR6wRIAWNmd6Z0r8+pPcz2u9YqocGa6IVIk0rZ5rMjf3YVXcnnQStFWiHnoJUZ/mrCGAISwmZczIxjtsBlVq+1ltHMHckoJK1nuTsaUOEyp3/lJQiAVPwZw1cynq2Osxw8+duV10a4TISurKqMrCMCd7JKkZsvZwqVJFFBMECI4Lw6V7Zd33P9bCbrZ90U7EUgYEx4ftaxXc54xs0wFMNeDwFJg+86nAvPc4WfE34+X8gLbtocwcy7YowtrW7myosqCnmmGGuICc/2nsXjvgEdbNvlWhdWbu3ff5cShk6SPRtIlDN2/c0v5+ZWI9AR6RiAgJ08fO905wEy5vglf25l7+MfXZzuXv2ZpsUHZBzdTO6d7/yBk5/XjBNaQKCC8csf/gcuIDu3OGwdf/xX/248GZAmznk2m4FkziAZIxGcVZY3v/J7/11hcYsQgXOwrOmob2eKldtffPB3f/b8wc80qRm3N7FtzhDByEMD4tKNN37lu/9D9favgJfzvEyGYfdk//Dl08ePP2yenyFqwZAjmQZRjowzFIwJwU1J3vcz19/+5tf+9f/EJEGo1cnZ6af33228uD9tN9utBiolirVMZcky7RyAr27uKzssbUw1XYdmy6cRGArLFUnp7fOuTzN6JWMlYyZm1UmcVdathHCV7tYr903/R8s4JETGLUSUcWRg6DQ+Qm45cAk9JZ6A0u5gLSUl2u+pnStJWs3cDCHwVD4Y4KqBGL0sdaVkeXlSEIACFHZGK2U72XyuAIgMkCUYffIubq6CwLXWCMkTGjtBImYmmQKh1gQw6F8QXG5kINKxnAaBjENMVYYxnWVUqS05uYoMQ+HltbA1QRyOG8/vG7F9KWOLiUpttdPvDnvns9TRiOwxhgzRcf2bX/wm2nnNbUKhtSYpn//sPw16F7brvvHV71jzqw9+9JeT8XAGI5on44wZZXK/WH37t75rZcqKpAYAy9WkG09+sXHvy7Wbb3e65x9870+jcAxaC9MOQPr04ECT5oxZnAsEvzT39u/8q7mN18nOci8bh5N+Y08wa+nL33r54Ocf//R7QTAmrSDddQyZ8ScW55bgDCFXqHzxd/6bu9/+Q237417L5YKi4Gh/58nTTx6/eBQEUwBQWgFqxoAxsDizOBecWYLblnAdUSxV+LXvfPfR409a+0/kaBBJGY6GNhOl2vLX/tm//Oa9a3NZ+8r5+Mr2mB3hhjlras4GajCRjzULzF49el/d3wlsxS0LAEipWfEBAM0Ks8jj1aN/VsEIgYBziwthHFF6OUBSAreugOmffQwZR8hFUiZHBAAToSUTBwEZw0s5rFcXMA23pkHFwBamTVfGMQD98V/+QKEtJ+PKwnJteT2bzdrCsgSb9fqfnbfO2m3PdhzPLZWKrmMDQBjH3U67dd5SKuKWkCgKheJkMkZmr27eEEiWJYbjsNVq2LZ90WtnHbs6X2Oz0JNAEw26nU7nYjruCSejAVQcIul4Op7fuhdMxqd7z+dqi65jj4Jg0msub9xIGkQBkkoPQRhHvWZjKmk6GSApJA1CEOkonNbWbnCtcuX5k/1n02FvafMGZwgMMBmrlv6mELxcniS1jnYAEW0HLUep+KJ5tPX21y2v0Dreuzg7WFy7nqjQMpbJ5Y0IJRCZqFEIp7K83R2OpIxIRXEwHPcubLTmb9xrHr9s7D2dKJibr3EAxoAZI2eYWAsyRBSMlRdWs+Wlfr8XTfpycO65fhRF/dGg022jEMd7O8fN0/lqjacdEIkOROoSOatvsekItFJSh5ORkynMr229/Y1/4vneG/VCJWOn7wtp+pB0dkgptVam2xaIEMAgs+YoEbYzy7P/C+YRxzGpmAkBRIY1mH4XMi6S1Bw/a2JEaWUwCgkITABPpK9iuyZPSGYVsM8xDwBTxzRYiFYKTBFEq1lxHy/DXUyriDMLTaIpw8gzpR6ttVbSkHz/3Q8+INsPg1GpXO02T5hU+VLJsi2bMw2kSD988ng8DYr5bBzFiwuLvuMEcfzzn/yo1+sdPX7fzZeICS0hXygMJ+NeYy/o9zu94fzCfCB1q3WWK5bOOx2IgvX1DTNmSAMQwUWzMe53gjCOwvF42BN+ToYT1CTD6bB1QCiiIHBsO1+oTKL49MWD1Wu3PTdjtjYD0IBxHB0+fbS6db3x7P5gMiIVAwAKgYxNeu2L3Ye9US+XLzuF0uHTj9xsvlxbNhjDJXgCSECnu8/BdpfWbzUOXwBqMAh6GLaP9ybHL0S5Ouy0L86O6utbQticXSZTg8FAa23ZVhhOnz/46PoXvrG8ebtzdhJPBjoOx/22CiNP2J3nH7cvTgInWymVLc7TZBgMLppUJQG63fOjvd07X/v2yvZrwXB4cfSCAVmWPQ6Ci+efDE6eds+OzkbjfKHkug7NAm4ENG2PW1/6rTiKB72u7WXufunXN+++02g2IZaVcuVePVf2bbjiOxLiCZCSUsmYlAKg5PBMJ5QL2+FCKCWvUoZe2d0z85CxlpHZfKTVFZSLWbbDhWUW+cwqiYERyDhK4WAgJc2gXbjyKSzHgLCIr0xfMwtopZSKGROccwOFaRUZhnwa5iESGeKjTmo+r8RTUsbIEqETrbXBqrWS5kX+7KefTKcxKlmeW8jnS3ff/OLJzvNMocAtizEWBtHOzkWTwwAAIABJREFUy5fAhe9Yjpcp53O2LT5892eB8Gk6aBy/yOSrwGAShhnLHo3601HH5ry4cffRh+972XwYK8/PToMoDiZzlTkvkzWodPvirNtqXrvzWhzHF83GsHfuetkwnKCOCNS03+nt3J/ffj0OAiG4m811eh05GS6tbbE0m1JKvXz0YGVzO5ct2JnM/rNPEQF1xBCBCIlUHMhBt7x63be8mPHjp/cXVjf9bA6S45cxJEn64OkjqWll82ZpYVEI++J4D5N8BbWMpIzj85NcfWPUu2g3T+sbN3nSsEmAzEiHBeHk8Scf12/cKRcKXjY/v3Z90G0H4y4HCCc97mds24kvTjuNgxGIbKHsON7sOE20ZBF7ndaLJw837r1dzGQymezixi2/MN/cfywnA9/zpePL8Sg82xudHZ4HkWZWoVAUyBEpESYg4OXbb8dhdP3NL9/94tdzxSJHLM/XDw9fBsP+r93bqvjJwMVLUR/SShquKzEmGOOJeQAyIZI5G8gMKeCV/PeKfWjT9BdHiWBukjlcIc9yU6fnZvLOzHWn1gHS0IqTioqaDdOc3cvEXeZhdEqwR5zlPhRHIUNzd0KWlH3Sj8u03LJd8z4qoSEnj2FaDo2egE6pzSnfDADw//q7d5vnLYsht+z55fXFer1UrR4/fWb5Hreti/ZFu9uTmvkWL1WqcTh98fDTs/5wvrag5bTROLaFrZWeTkaco4yCyajHuZUpL+Xm63uP75fnq9zxwjBSWmVdt1QpA+LF+Vnr4PDGvTeEEEyI46OD8eBCeDlOpOMQERjnJCwdTTbe/mb35MB1HWVljp5+tHHrddt2TPF35+H9+vpmvlAGBpl8edRu9UcDYAwYM5w6YFyjJq1qm7dBykkcNPdfrBh6ImOIKJXafXAfbWdt+6YQDIGVF1elhH67wYRgwmLCQmGj54XNw1x9fTroXrQa8yvrglsMGEMSDINo+uT+R6s3XisXijbnCGg5Tn3zzjQIx/0LZDwKJl5xrjC/OjnZ6RztdqRyc+V8xjeq2ybWajVPnj99cu3el/IZXzCOgFzw0vziwvZr/Xa72zzwhJ2t1kVpbnz4NOyfDaOoNxp5uZzveQKRIUgifvvb3733ld+Yr68yxjgwxoAjFIqVxsnp22ulerU44yYQgdJKSUlKApFhuc8KZ8KyksbUNA5NQpcUYro8vDVJGWkZc84NB/MSOEJm+q5moBMimw1oRkzSQiOnkN5Cwi+FUAwvZRZmi1zm6QBKxpq0SXIY51pLulL4T8yJKGXyJgmJvvI9SknzAEnexZgBDVILw//zb/+h1WpmMgXHdle2b5SLRVvwAOi9n/ygVKk2ztvTKJCRymYcN5N59NF7fmWhslCnMECQJwe7luMx5GEsfcfRSgbjHpC89dY3bMvJlefOXj5zPV9y1ul2S9l8ZW7uvNn46B9+duetL2UzHgKzXLtxcjyZTuIgsP2MDKeIZITp4jhaWL9dqq1cHO56uWxn0BOg5hdWAWjvyaO5haXK3BxLscdidWn30w+1bTOgBOfijDExHXZz1cWF5c1Bq9kbnMsoWly9ZvoUnj340PHzyxvXuUgpRQhzy+vDfm/UO0dkaBoAkDHLDZvH2aX1ce+i22vXljdsy0LE0Xjy+ONfrN24VyzkBWOG+sAYQ4a1teukcdg9A9JxMCZuFWsrwfnhsHXcCqbc8Yu5oiU4kW6eHO88e7p9762s71mzJlcDiLve4uYtZjmNwx0ZDDOZolddHh0+05OhQuh02oqxXDYPgE8+epf/zv/4bx3XQwQDDxtWsyVYqVJ7a71SySRKMJpISaWVmpmHiSkIABlaVnrqzyodZk8zliTxaWSfoF4yTsN3SksOgMiMKFa6Q81/wMRgJgkGMwDRlPm5oCvTzSH1dQgobHtGFzZ/MMZMnoOMaa1NAQQBhBCm+/dVB2ISXxKp5KZ5NWRoBswjYhzHjHOT0ptiCGlFSdsWILL/+0cftZqnxXKVCev6rXu+5zJk3f5Q2dlnDz4EIUKpAZjjsJPnjysLq/lKlXGxtrw06nXOjvc8x+eWNZUq5/kaaDoeopar199Ebtk2d/zC4YuHruf3RpPlpXoUjO+/9/Pq+vXqXMX3XPPKg9FoMuz1OmdevhjGE0Y66TKTkjtOZWkzX6qc7jxm2Xzz5dO1m/dePLyfyebqyytCsJQ9ymzHlVF03jjggiNREsUQIcDgorG4fbdQKDWP97qtk2y15nq5px/+wi9W62vrtjCpcpr1Mja/snl+ehJM+sk/Mk4cUYhp4zC7uj1sngwHvVp9rd8fPLz//vrN10vFvCOE0XNEnPHYca6+ZjmZztkREak4iEkXaqvh2VHca16MRgFgvlBqHOzuPn+2/fo7ed9PZ8qYymRyWHPGKgvLtZWtduOoe35k2Va+ujg62tHhGIU97HUGo1Hz7CQIJf/qd/8NZ4bxj4IxDmglfUD4xnKp5AnSisDQY5VpJGTcgmT4MDA+IzulmfzVOAXR1NS0UsjQRGiU8Pw40ZVj2zTBG2T5SiUxdQKo0wGiMo6AKDGPhAl/NVFCo981czozp2YiJa2UUpKAGKCwbEBT/ZgBxGmsRsS4EMK6iuSZpQxEQUQIBEbW2lRGlDL+xDzxn37/vc55a35123a8res3bUtYnMdI0zByvMLL5w8G3VamWGnsPKwurZfnF7gQmiCb8Qb9zsnJfiZbtP1Mf9AtFkuIMBn3lYqXtm4x4Vic28JyMsW9J78Yx7EOhvvPny2u3/J83/PcQsZPKNUE7YuLQfeCMWCCoYrNcU6IwWiwdP2eZTleJrf/4L2IdOtoR6G9sLRSKuRn845JEwKUF+r7D96XJFMCYBJp6jgajQert992Le/s5cOL1unZ8Wl1dWtlZc2xLeTIMDn8zM+Nc7GwutXc3w2DMQIiaQYIwBjn4+Pd/NrNfuPo7HjvaO/5tde+VK3MWcJ4rHRnMeA8IekWqwvZQqXd2JfxREWRiqXlZ8PWsZ6OBpPx+WAw6HZu3Hs7n81aliU440kf1VUoAQDAzWbr23e0VOdHL6ModBwvaJ2oaMocPw4DqVW2UmWCo2BgMRSIHMn8VXBmCWQcGeeaQKk4ofGRNoOgTbpsaLafm5Ff/buhuEspVRyTkpDMub00D0ObRZYiTlcNLTUVxjlBMheKcW5ws+SFL69AnkK3n30eRADgnBvECYElQ5yVJqVTv3FpI5AMdoNfejNgjGutAZEIeFJIMSR/lVopAEE0GSKpcDJUSprRi4iEmgTjrufUN++Mp+Ner5XJFUtz87MBiK12L45DHQXjcW806Og46HVbk2EflRSkZBgkQS8jz7NWb7yJpHfe//5cfd3zHItjHEtkwBhjyMrlynQyYqDUeMiVBiUZaa6IKx0P2p3DpwiYK5Zrm7fQyQ3Ojuv1VSmlVIqzpEHPAIGO7b75jd+mIAZSKCOUESOFSqGUnRcPdj/56cLW9cWbXwzjeHz8eK5UNuUrw7NjiDytXjNEP1P46ne+67sZkhEoBTJCGepoCtNR95OflNa2h5329OgJV6FgIBIbo9SLmLIPmResb93+0m/9V65fpnAaDdvjzhkCwaAdDzqj1jEJiOLAtYXFCSEtHyMYU0lLhAwILMu6++VvvfPtP7Dd3LjbAiA16k+n0yicxJP+oLGbxpaIFmMiFVdGJKm1GZsGpIGMWreBWDVphYBCzIhSn7WN9Mx99Z+SLFuDIc+ms5gRmTAdJr8EyM4+khsrCQnznEhLY6aUfpgwLKGHfM5CSeCglUy9ASciJU2FkQBmj2QAFZamQ5cvYe52+S5X4jjzAOmtCACC6RAQxsMeAAmWkIIjqRiC4OhYHJQMRiNJmgvGePLMrmsLZCQlSRlHESHGYaClZKRBqXgyovRFOBeoZDQdIufh4ML0gcdRRIQGX/M9J5vNZ7P5MJwwy+HcIkBKnf/Bww+UlkRaadLhMIyDcfeMAUyCKYOkeZUxMmWF5Ru35xfXkGzgqAEN1VqRIlAHH/x963Q/iiQOB+NO8/kHf8vMdiFiYBRrEiqEqfpny5V3vvX7tpMHLjQXxITpL9BxOO02N7/4jZjgg7/6k9GwA6CTaX2kOSJPafOMoVEqKy0sf+Wf/2GhtkVMMIbEOAi7VF3ktn/RONp58tH+0S4DSBqHEcwYh6QEwcAU0Rkggp5f3vjK7/63K1/8J+gWgItMtjCehKNeVwYB/9V/+W9EYltosGSp1TgIn+0+f72WqZcSDbKZBQMgM9LujP9jruMVKjuQUsrwUBDRoF6AAMAAkXEuTL/4LxcsruzspClKK/Pj0TJOF8ErRYsrkg6vOrHZh5JSJzQqI06lTGsHAACwJP1gCESXROAr72UsIelDvOyiZgB0hSpvom7+J3/+PVGolWtLi8sbS/VFgYwhNLuDWMZKxS9fvgiCsDS3qJUUnGcyWcY5aaqWCqdnx81Ws1hZzObLkyjOZDKu6wdhGMdhcW4xW1rgjAHiZDg8PtnP5io8U5CTnvAymWyOAH3P8WxbAzBkkygc9HrD/jn3S2auiWkLJaBw1M/MLzYarYX5mq2ikdTd05d2ruh42UI+J1jCYjTbW6DIVxZ2Hn0InIM2uSMBgY5jiKNh++zGl34znvSH02mveZyZm5+rLlJKE0iOf6DEWAgyhWImVz54+VDFoQpDHU6IIVn2NAg9P1u7/Xb7eO9g58nq9i3XdRGZ8diGz4SMIREaZB/Icf3FrZv984t+6wSB0LYn03E2U4i5NRkPp+NhdzpemKvatpWyPSB1SMnbGXMhAibshY0bhZXrnV6n3zq0LTtUMJkO+W/84R+ZnjfGEIEirc97nQ8/+cXF0e63v3BrsVJMj85EOYFbdiJD+OoexM8xDzL5/Yz8k+whTBLqhAyffnzelk7OZdNngoxzYZFSkBzk5gBPKpqJ9sI/uhAQaRlFwJgQJhKjhH91eUWSoCMyMzP6qnkYP2akgs0wADNy0WgIaSXTSigCY4DwJ3/x1yxTQWatrKzNlSuO4EC61RtKGR0e7AkuFBe+l12sLgyGAyLwM1nSUMx4ne5F4/TY97PcsqdB4FjCFmIaTnU4zeRLucoSF3w6HjUbJ/WFJWQo3KyQsbDdyXSay+cJsZTLmsOMC/tgbyecDrVSwnaVClOlAa2jSMl46+47xWwuk8k1z5s6GJbnl3u9nudnc7msqZeZI4iA/Fx+0utedM4twTWQaTbQcYyIcTjljrd570u983Pwc62Xj+vbd3wvS0TGdQBi0jhlYFiCYqXGuH26/4JkCIhoOWi7ADQdjXw/N3f99fOjlyeHeyub12zbvZyzeqX0m+wZAsHt+tadIJLtTotbFkc+HfU9y82WqpNgGo76rUG/VKpkPE/rdFgzaCBkiIQwo4+bmDBXrNSvv0YKOicvVTi23JxpcAdEiJWaxPLx7ot33/1RdHGatRJq8Mw8kDHLTnhW/5htzMqBhnmopDKlQAQwUKlxVCZTt4xk8ucf94lhGvNIJuJaVlKjZAyu8BwIjfCu+LzgamYgIOOYEExDAZjnIXrlm9Jo8HOWQgAgpbUmDUCXKA0mAF0KBOPMorhmRo8+XyzKMBQcHc4J9Onxke942VzOlIBtWywtLo8m49Z5S6pIMCIARgpVzLXiSEppJOTIJIMwGMYy7LbOTo73l5fqruv6niccN5RRsVjiDE9OjybTQGnFETUARSEXlp8tR9MJMoFgE3ACRoSE0Dndl+FkEoRuNlcpzkGmNLo4KZdKT549PWmcIrKrkQVpVVxYgVgpFEigpJZKo7DAcsFyj5/+Yjzqv/GVb5Wq9VDRRz/8yyiOZhyEJNQxBpM29tx686vl6hIwDrbHvYxwPGHZUTg42fkk6pzd+JVvTYPJz7//vUbj2Ayu0gY2ZIhAhjyW0hzRsq23vvV7K7fe4m4BuIVIo85x73jXsW0QVqdxeP/jn+83Tgj0zvOnrfYFpCQ0nlgIcI624BbnFuP5TP6d3/idt7/9+162FIdj/vrv/uuHz54Vi6VRMP75x79oHjzzSTlcuF7+q7c3F0q55Kw2eqRXdHeSHfWZgIZIaW28hxmKgMzMd1WX34Om11Wkwor/JfNQpvKNzBS2L/P7K+lOqoDB/7HFjLhjIq+aOuyE334FqJpZOhpwMEWKjb8iIqU1ApIm5CwheiiZRFkqjR4xaYn5P/7mhzxTIaUy2fwnH/zDyvoWE/z+pw8dYWWzmSAKW80TrnV1rsq5yGbznV53/9GH40nQazeH47HvZ4XjTCIlEC2bh1EUBFPOkHMRSSV755XFVfPb7Y5GQb9dqy16vg/I2p3O0kLNsa2DnWc/+MHf6mjCPH/cbohsUZHSpBVpUgoQiGA67jdODlUwLc/VBtNg0D6tLa2WCuXTs7PecFApV4TgiKBI737yUXV5ud04Ggy7iBxkTKgZNyKsgAjd1ml2bkHG8VSqfuuUMZyvr3LOIOHZJdUIk28S0M6nH1S37ggQw26LGWskQK1lFIx6HU5YriycPH7/Zac7v7Se81xkzKSapkNhFnoY2nXz9DCK9O0v/lrn7CgORqilDKfBoOtZfr6yOOyejzoXD3/0nxTJJzvPCnO1nJ9J9H6IODIwesHGIQBopV4+eXD9y7+5ce0eb2bnxp3m/rNPGq2mGrazgruuj9w9P9r99bduLc/Pmfje+KCrLa+fH+gTxXFk5AmNxZvfCFzuNTRjN5S67D38nAUJwExtj2MAwjRVv/rNxj5N9cPULj8/WiNSWqk4Nl9inGslSSm6jAcvkWkjimc5rlIqYfmkGbpSmpnyZYrnm6ZCMuNwjZfB5ItE9Kc//IUkPjh+LsOpzs43D54NIh1FcT5XIKJgOp3G2vf8Qr6AnAHgoNskrTnqnXf/k52vCMvl3JqEIUducZQyDoNJNLjoPftoYesWMSeeDP18kQGEsZoE41I+b1mOZTuA7KLdtgR/92c/ntu45cRTBWw8GmhEy/E0EWgNWiEwZDzsXdCg69e3mI5t2xmFkcNUrlj1PD8Mo8k0rFbKSHhxdhrF0ermdT9b2HnwPvOyQBIAGRfITVMJoyho7jyYnB/n61tS6Yvj3dL8Uq5QNNOzroRGBABnR/ujyejmrTfrG9udZnM86hnACwCRSMkoiiOmwqjblP3zPtjzi0uuZTFkSQWOzTYAAsKo33/24MPX3vnGXKW6uHm73WpE0zEyBNJhOAElC7X1OAp6Z/vT9oml46OLjpvJ57IZk5Yk5VGTyyJorZ99+gunWFtf25yrVLhfW7VBX7x8WK0t+I5bKFY7zUb37CCcDL/z1XdWlxYt22EJi0SmWk+/hFMlGbmO4whUbLqREFEbrm7KjwbTx2s7iMg4V1KydEW8msCkIJWUMZhOjyuMxgSqSo4k5MIy/bEJM+qzRkKmBqKJjH8nUmToMHC5jLFcBAIiYdtGNkZJyThDMzRdKbOsUjLpFjHIowHH0t9Y4s+Qkdb/788fExOZwsLi9m3gdvO82b1o1VfWEVBrNZmOQ02+bedzOUAcjwdnB8+Xr72mVNQeDD0/7zquZbtBHAFCxrJJx0EcSi0BFAe2fOed1uHzTC5nWU4YRVJrG8nzc8CYJZxIy599/z/Pr9zIZnJzi4vDi1ak1bTfyRYqjICUNNPrkSMyplVcXbsuCAvFwjCMe2cHtfqGkV/iQhSL+eFk/OO/++vX3v5KznMzhXKv022fHQovg6QgqeLxxBVzHo96QaeRX9mKplFr73G5vpHL5ihRRk6O/36nvfvs8d23vuJalhDW4taN5t5uMOlDcuQBMKbjQCEvVhbDQXt08rJnZaqVeUvwJPcDnbYXUhhGH/3Dj7Ze/1I5n7ct7nhOffu1fq877p0DkFZxHEwhHDvZfK6+OTw7lr1WMGyPYhUpKJVKFhfImMG1ibTWtL/zpDea3LjzuucIjsjnbr4+PNu/9oWvloplQNE62Q8GnSicCNv/nd/85srCPKZwHWNMSslnB/8s/AAAICmVUpKUZMi4GalsCCmvmIdBrhL0DxlqJdmrnsQk50YxhJQ0AzH/sVAMGTdToMxx8st0SZNPKikxrfeTUlc94WwlRCStZ5UZRDDiq5xzndqnJiKdqJVqrbkQphXk6gMZCgIR/dUHT2LiwhJz80tRHLvZXPtk3/N8x/WUptF0Kgl92/Y9V2u99+ij5Wuv2Y6vdTRsn2VyBc/POn4miiOttOc5iJYkqeIYubBz5aX1G7lC+fj5p8W5BaWVIq7DcT5fAs400OHOw0yxWixXCaBcLg26beRW9+I0X1rwPFdqTaCBM8YF4wy4JeP4xhe/fr7/XLh+fzLJObabLXDGiTQhvPeD70V+MZ/NVyslRCzX6k8++UC4nuACERi3mBDIODDkyLXtqPEQZJCt1SfBZNQ+X9m6bSQMze4Po/DBez+9+/bXshkfOSAwi9vV9WtnR3txHDBumSoMIMo4YF42V56fnB30zg7GfqFWmReC8aRwyBBAkf74Zz8s1DcXF5cEZ8g4IAguFjZvKuK95qkJPaI4YKBB6dzKjUmnGZ0dRFpGhMPJpFgs+a6TZP0IjZOT588f3XnzK1nPsQXnDLmVL9z50q/6hXK71Qomg8mwK+MwP1f/ym//wdfvblcy9isbAFAqyVKhqhSah5l5IKJIzWPG4UvMwwzFTD2G2bAEYHKVK5saCEBpqWSUnNP4yxvabGojKpd+FYHhpV9KbQ2UTFAmxjklqcjsVslLYYplc8viiU4F6BlEkdqcobUbWzJtITONopmZIaLB/v6/nz+eRLHNLb9YimMlGHOyhf0nH5aqi4zz4WikAH3bdl3n8MXjbKlaqtSISEfBRevENvuP80hqGUvH5oiglYzDKSPNGFvZvG1xGxB6reNscW4wCeNJv1KZJ4ats+PRcLS0ummmQPpeNhoPwigYDvtA5GWyURRKGSGRAOSAgBQH47n61tz80tnLpyyTG7Yb9foGMk4Iz5/cb/WHtYVVpXRtrmwL4XguINt79LFXLIPSQJqQEI32jEYEbdlRu+mXq4BMhgFjOLewjIgMmdL6yS/erV+7PV+ppHoggAi2484trZ8c7CoZAAAZ7IswnI4sP+/6uenp/qDfGTu5pflF0zqLDIno2aefxGhtXbvtWolWGQMTDrBqfc3NlS9O90mFoGQwDWzBOWjMzoWDc9VpMtcH0t1B33G9fC5HRO12+/57P7n9xW8UszkueFJbfPM7fxCRiKdTFU2HnRYQbb3+1de/9m0vm399KV/2rVkYkgYwqLXizDSdgyZQSiatS6SZsNKgiC6NA4ALYVmXrSZwZcEE4zI1WCKaMa/0K6zHXzYQU5O5ar3GL82MhNJEHwzF0ARsn+OOTFmKzJoJ8G7KBoAJQ5mlIRZnZCQOGNJnO1JSBJIIAP79D9/vD0aWsNxCWUklGLcYJ2GdvXxcqi31hwNmuTlHDAf9Yb9d37hhNIRkND0/PRDC4YjAhFQyiiKXMdQUxVEUTJCUJr28dVcw5mcL7dNDxgXYfjgZVCvzo9Fg/9nj1Wt3HdsoWTLLEgi6d3EeazUcdPP5MgApGSFJ07JLgAikCNavvx6Nh53WSQhYyOWz+WKv33nx6P7i+g3P9TiiZYmFUt4TOD9ff/Hs8Wg08HN5hmR6+5ALUz9njIPrT072KtfuTdstKVWhXM3l8lLphx+/HxLcuH7btni6BUy5nbxMplSuNU8PkHFuWUJYTHDkPA6n+doKIzVtvBxOplMnU6/O2ZZQUjcbx4f7+7e+8OWMKxIp6/SMMrupMr9Uqq1cNBuxChEgCCaCi+r84lhRdHEqx32WKzCCXq+nkBHgez/4641bX6hW522Li5Snwm9+81+4uey0ex4F42xp/s5Xvr12+w3XdRlj95ZyZc+6/P2ne8A03iIykyqY5iHQKpFjSwKvy4SBW5ciKVe3Z7IgY0rGiGj4FEprrSQYxi4zjauXwMUsb+CWlTT3vbIaAaHSirRijJsWwuSpGTeyiwifZyGIoDW3LGGmXgCoVNwecQZYgVFwREAzQD05F9Kbz57T+M7/8KMPh+NpJpe3MgUgZXo7hWUP+t1+90Ih95xsHI1Pdh9u3nnL9z3GhNIUBcPzox2LCfNTDoNJFIacYtJaxqGcjrQMKZZLm7csyxUcM7nC/uOPnXw5DCae5z998F5t/Xo+mxPpD1xpnfXcxu4z0vFk0BHMFqBVOKU4JC1JS1CKlJoMeotbdxbr662XT8dayuEgPzf/6Xs/Kiyu+67vOjbnbDINNpZqnDNA4eUKT+6/xxlH0KQkKIUETBNqjYaYIHjQOi5t3+0cvAiicL6+trPz/P7H783VtxcXqq4QyQYBAECBnAByxZKw3ObRLigFSMaNAOhg1HWrdTXuRxfHvTCccK8+N3fWbP3i3Z/c/vI3y1nftkxWAiwNHRCBI0OAXKFUqS31O504mCBSFE6H4+HixnVmOZPTlzIMrGwBGYwHg7PzViZfXl3ZsG0rlVFBxpAvvf4r/eahiqJ8tX7tra8vrG5wxizBEeHuQrbkW5+tDCIiopKKEjxXE5gJByhsO+HqXsFOedoqeAkL/xJoZdpFjL6OUjEpaYIrTFS0LgUOzZ416hBXbWNmfCZfn80Z1VoDEBdCq/hKfHf1M4maANGybUwkQ9OG+9TBKCnJ+B8iYVnmmNBaJlJ3V52syWcY+/N3P51GcWl+CYWFYKRAmOCcO/7JzsPBdJItVI4e/EN9+7VSuZIOo8MoGLVO9h3bNUlCFEeTydC1HcYYKRlHgVaSSM4vb7l+jjN0LVsRHbz41MqV9j/9iV9cnK/VbcuGZAQ500oTsH7rRJEOxgOlpe84ZqaKqb2iJtCKZMj9XHVpvVgs733y8+F0dHF2qCxvcXHN5sxxXYZMabIsq5DNaIJ8qdw6PW2evhSMMU1GniYJH4iQNBJGwRiROZWl9v7TVuvsyacf1rbvZWxHMF4s5lNxjBQLRkDd/foBAAAWk0lEQVTA8tx8HIWt4z1QhlWkkYgRxdOx5efjXotGvZGigYSPf/S9bG11pb6Wy/iCYyJ2AkiG9mHSHoZA2s8VqgvLneZJNBmSliSjcffcyZfloBcPOxK07WU55xaC7WfcbC6b8QTngnNTK+S55TWpVH5p661f++1CZU4kdwLG2J1aJlG2ntUMrhiK1kkInlbx+CwtmX2TKfO94j1+6QQ3o220kU8nImW0ToBzjles4uoutOyZdNUVMCrlZyXLKmlQZsZFQri6ioMlnwySmErNHAiYEOuKeYCZ0qaVES4zzfdgKiqXhj9zcQCkkfE/++nHoyCcX1qR2nCckDNkgDZnEbcv9h/nFlaDQWd165Zj22YRIoijyUXjgFsWcdAMNempUo4tGEPQKtax1hK0riysZIpVzpAjCNs5ON7n2cK0sbd65+2cl2GMQ1LTBEQWKslADgedKJrG05FdqlIcxiqiFEYHINA06bfr1+8WC8VpGI8ZHx89q22+Vi3PuZ6L6Zk3mk5rlbJtcQIo15afffBjsD2GBFoSaAQCTaiV8U46jsKz/dz6TcqUB/tPBNLSxi3f87VWwrEyrjf7ieEl8ZbVltfCILg42jUwOkmpZaziIB4NdDhhcaSkHGsqLSw5lucIK+t7vudeSqOniMwlhg/geP7K9q3uWWPYOoF4CmEw6TTiUR+00lKRV+CCccF1HEwmY27ZhVyeYdLszivX37z3q//87pd/1bEdYzVJvyXC3doV7fdLOJbMBDPjAJL4yvycMSHsQML8FcKy4DNH95Vjn5IGEwAAIkpaOK50KaUsPZrRHAHAsiyeph9X4zaT9Ke7mkhKAjTpoJaxaWkgurJUsjYBaTSc+TS5UpdacnAlR09ymCTJMdHgjEiA6WuQNpSmP/6zP28c7S+uXiNmzcitQBSG07Pjl73T3YkCNen6pVrG93kyHVzHk0Fj96GUMgyjyXQ6mYyBCy0jGUziYIhxxEkzoFypWqzWQVNv2H/58mn3dHckGXWO7ELVsW3T6EtpaBpJiSCP915EgzZOh8wvgoyZiphSjMiUyTiAHA/dYuW83Ts+2pmO+nrYIxUBsxM6DzNJI0qtq+Ui+//LupImOa7jnPmW2qv3ZRYMMCAIkCAskRRFyVs4TFrh8EEX/wDJEfbZpk8++GfY/8AHhx0+MEIORShCJmVZFLSSIAkJBEmsBGYw3T3TS3VX1/pe+vCqembIOXTMYaaqujvzZeaXX34J6HpeltMXd2/Z7eFpjYeoiyxfRSpZQZ6hUvHJaPjS6/PZtDz8zGt2g86Ac15kme8HtpSb6GHQSDNYtbV3ZRpFs+MjQoKq/CaVxlBkBGCFXfDbwnGFYI7FQZPlWK5dTcUQwWbcdHNZAOBc7F17KS9hfnSgodRFQVlCRMilDrsamWRMcMG0iqMoLop2s+lYAgH5X//zv2zt7XPD5qwPQUTgDG5s+S1Xnj3+TWdAV0SSmqtbY1a4SS0RhbA2C+bO+cbG7Kgi0WnStSopIeDprB9CXTWc/jMXsiKln3cPINA1KGu0iQx3CxGBNJCuAshZB908LmnkvAIS0EBY1YpZqLQdSOuqd47IDLtnQ7/fdFVqIAsAgHH+w/c/RzscXHquKEtEIK2jaDYeH43HR0WyTArqXXwpX4y0sMfHx2meWbbDuUizeDwZhZ3tsNkLmh3H9TMF/d5Wszu0grbiMteqJG15oXSbjx5+Fi8XzbC5GB809q5l80lzsBOvlsez43gdE5BVbYRk0nEdL2xsXT5ZRrbX2H3+ReE2c2HlXCghNZeKsQIpW0zbF666trc6uF9YrlUm25dfTJNkHs2i5XKdrAl0VqhWq+naFiE1+tu/v/1BUZbh1gWNjIQEIcmywfVIOqQKIq2RNS690BrsLI5H0cHn4Pgm/StK1Ww1+Znyuv74kBCGF55brNZ5kTPHA9spGSuzBEpFjHn7L1278Y0Hn9xy/bC0rPjkuMgyaduu6yBWTW2sRlNq96szua2959zO9tH4SOlCpWsGQI3O5RuvL6fTJIkd1zWslmwdzeO17Xu+4/A3/+6fOMNaZ6LCARiiQHxpGJx6CIEmUqqsGnPmwEYwCtPmYeo3y4S0DLXpy7X5aWgwaqBaaw0Epug3muq0GWaqobNTmMrsVq/d8Zx7kDbGXNdFJSFDQM55rZ648ZBzCZsJUIZQYy5mpoLNE1KtU6GVRsYBSErLAGhKnR1LrN3+tFPE/vN/fpHk1Nrenc3nJ8eT+exEcN5udbqNFmm1TPNmsysgv3L15Warwzg7OhofTY5sKI4ffYZlptJ1ma6y1bwgknkCWZrHUbqcFeuFzjOuaffa11qNTr/bbQSN1XwiHB+I+t3uYOtiEDZt241Wi9FkvIrjPM9LVa4OH8Tzk2w1y9KYSp2tFvlyqpKYsjUUGeQZZGm+OLl4/dVWs0NlvkjXKom7g+3BcMf3Q9fzhZRpsj6eHj95dpTlebvVcl1XuuGnH93UZYlFqrK1zhIqcsrzMltTkSOXXMgiS698/dul5a2OR4XWW7uX1qvVaHy0ztJetyurFhszlR4BIpIUsr914dFnd5LlVJe5TlPKUkIg28qzjHErCFsnx0cMyG40OcHxZJSkKRdCWpY4lXg7LTgNmQiBNzo92wsPHt5TRcb8BtrOMl4NdvatRn8ynfjSQoYcWZnG00UEXPA3vveW4AyZiaLACaqSB6DyEHNiEpVluTlciaomhq4xn9pMkHMpNu5x/pgHIK1JaaWVpnrlNiAYPaGqRXWql1VhWXWywGQ9W3sOsK321qqKL4xMl6XJh5gQdGYIflMSmqthnSwhFxtFLF2NChLCxuE3eLQZTOBVaFHqTGHDwAAfjJFZq8v4Dz98IPzGOi/iVdzvdPvdbsP3JeeIEMfLNbM8x7cY9QYXbFu6jtdsdYKgoXU+mjxzw7ZwA255CnmulB+EtuMWBLku8zID0pro4vVXbC4tKTnDrChyYpbjY5E2213OhW1ZQdBoNpqu6yqlirJsBl40n5Zlma3mfmdQlrkqM62M6oACrajISBUg+ODSC5a0o/kM/YaajTu7+2anMePC8/xWo+nYzny5aoRBKwyaveH44OnseMyEoDzVqtRlSWVBRQ5Gu4zxQus8mu2+8AdJSdHTe7Zl9bYutpqt2SL67P79dZoGvm9VGVdVjQCA5TjDnf0Hv38/jWYqS6AsAJChAF0W0UyXJZYFSjfPU7CcVqOlVXkyOjo5mSkiy3Zswes8p2YW1vG+0el3t/fGj+8XRcqIKF1Fx4fraGpzy+kMOaAqcyEEFVkUzfkb33+rzowQDe0WK8Lti8Og6QjSVCqtK+GfTb6tDVZk7r+xWCGkKc2/mlxp0uUZO0aj1m4S9yobUnS+fX7Wx4SQtbrcmYfQVKqStGE0ICJTWlcZEeOMcdqMf5x9rQOUwWqFsATnBFQUpda6HtM5pfcrXRoyIucCa8H5as/o5pOrv11dSVyzH3382PJC2wsC13Mty1BVGKAmFa/jjNuhG0jOmq0OInIhTNQC0Ito1eltB62eFTSF40fr9WC4E7Z6XtjUjKdKI5cFE3v71yQTUnDBEJDNo4XfHWSLSbu3xRk3KhmcMyGkYzu27bZ7/TTLWdBYTCdO2A47/ZIJjaiQaQNXEAHjaZJcvP4yKN0IwsU6W65mg/5ASBcABecMgHMuuJRSpnmx3e9Kzhv93Tvv/1yEbeb4jAtiTBkAhnGQFtg2MAbScaVobu3HSscno0ajYftN13Y8z0/WySf37rme22w2wMxeARhYyvb83t7VR188KPIYkINlo+UAl8RIMyto95P5VDEhUHMv9C0nDEMiPZvND8eTQb8rhDhtCgMgImHVgPbD9oXrr0zGo3w1RzTz4QUXnNbLtNSNTl8VGSIiKf5n3/v76qgko/oKZsEhMrw+8EMLTRq+OYXpbJq+sVdERJSWLaSs0adzx7yJQhWvzwBPdVGPYEYO9bkxvc21EQCAceN459yjVJVHbXi4BjU2aS7nTJcFfeWCZ58JNAGitK2ak0WbuLG5jyatlWKCY2X6ABUvmE6vA2QSUTh9C/Tv//1OQSCcEBE4QzPIiQQcYDw5UsyygVzH9sOGYRwTaK2pSOPjp/c5AOU5lYXOk2SdOBy51jrPVLoukrVWBRRqsHvJclzDAM/zdDJ+Jr1GdHywvXsRgBniBlU9QSAgyVm2WgnGknUcJ1G31eWMkSpBa9JKqRIQ0bKBC78zsN1QICPEVZarPB30t5Fz0lpwAaZxhawoSimtVhjYnrdOisef3/aaXRBSISuU1siE6wnPl7bPhFS6KJi1fel5yw+Wi5lww053IKUgAMF54Id5UbTbbVmrp2/OnaARMm49GR2S7ThBS3qBcF20bEUqK7Ptqzf6w72jo8e6yMj2HNtq+KHtuVrpLMvDMOSM1alyVY5oIEQQjNmOs/f8dbKCtCjRsrhtKwBwguH2pVITN/ohAPzNv/lHqGEE07+O1itCyLLsWtfteHa1JKCya0MIqE7hTQIEde2Bp9DVeffQlcynGQHFuq22IeRS7T9nj+RKN4+d5lenyJXpu1SpJhAQAiiliIAzXs3p0AbOqRs0VUaEiNygWFxaxsf0pgFy/seQebHamlu9hTOt9NPCY1Pcm/v9x7u/BLc5O5lwxmzbFowxIxmj9dHRF9JrY1najvS9ABCJYHT4OEuTPFlNntwnVRTpOktWebzMSwXpOlvNktUiWc3SeFGmMeXrMGzHcbqejZq9/nq1ihYzp9FbjB/3htuWZRMBma3ZQLPF9NmnH9tB4+SLT6PjZ/l6mccREZSLkzyeZ+tIrVdYpEIprkssiziKnHZ3vpgeHX7R39kfP7jTGmw7jiuk1KShNgACWCf5sNf58Nc3jxfR6vB+mueULFWypCzBMmdaY1lCmVGRQZZli+P50cFw73kunZOn959Gq6Yf+rbFOFOalFJ5nndaLSODvJkGKcviwce3fK+5fPIZ5ClliU5jShPMUkqixehptpj6jR4yNp+dFIyjVsky+vnNn/jdAWjtea6sOxtQdUuqgoIhWpadLeeFBsgylaxB5UWynB0fqrIMutvS9VWe8je+/5aB1c3JGafZ2+/8+ODu71aL+bdfvDQIHdgEhXrN2vmmBwAg44IBshot/dJprTXRhuFY1TOVOLwRdKOKlgvnMpb6hTFuOgwbfzBJ3hmclxDQGB8gGmXUKifczDlVoAbDWsjd6NBxxkulGMMzk+enoQEQDA3egG+m309aY61TYOIVGjYd48aAjFbMO/dPPv3Nz+zu8OjBna2di4IxJEQAlReT6cRpb5PKHcvy/BAQ0zx7dOdDInXwu5vh3out/q7fHQadoWy0ojzrdLfD7sBrd7nbyIVV2C5azvzB74BDFC2GW7uqLNdJbLmNJFl1W20mLASmzaet9cM7vw2He+vD+8vjZ+2d59ALFtNx2NsLOx3FZYFQAgMhmGUzy0HLLopsevumVoUzvJxOn1ntgYomveEFrCsEqo4e0FrP49Uvb74b7jwfoj4+fGD1LhQqJ1JgkjzOkTNCJAZAoABYlp7cu6VIZet5a/eKK6SZrGGcpVmOjDWDAIAREgIQ4MPbt9o7e6+89u3RyTReL1BI4JxxDqwaiSAAV1jL+UR6ASTrz3/6g+H+c8nJ4WidOm7AAH3fF8Yyq7IRDbsUGebx8vb7v/6jv/jutRuvTI4OlqOnVBSUJ0UcpfPj+ejQaff5d77/DxVUD/BsOnvnF+8dvv+/bd+9/e7b3/3zP9nbHlaxybTPv5K0MMYt22GclaXacOPPBpDKPcx5TKSUQq2oWmeDxuBqFYUaO66UGQCATGGjla6waERzTaBTc0ZAIlJlCQY20GXd96i7iOcaIJWLAREyxqXRYSm+QjE2GBYpXZqR3apGMgX6mQwLN+cF1X8DAED/9c5NrzV0O8PJ4UPPDbwgQETShAwORs+CznaxXjYaoW07GvXDT293ty8BYKKoETRdx7WElEIKIZartctZw/MsLoVBAgiAlLYsm/Nw53J09KTR7pVlqYFpIptjEDaUrijS0+loNj648NxLveFe0O4L23O8xiJZ51nWH17gllNoUEBCWtx2uXSYlMgl2XZ6cL996UWVxNIPy7Lsdnq24yilNIHZuISImujWr/+PBe1hf6e3d3l89HS9XjWG+8J2uOsx15deKJyAOT46DrNdEqKw5HBnf/bJby3XXyrV7g49WwKwUmtkLEkS1/McxzKQbRTN7t298/I3/zDwnL39K8fTqCCyvMByG8IPuBswxyeGSsj9G68FQWt0PKJkObl3e+/6Nw7u3ircJkgLiqIRBoKzqrlS4zVa0/vvvXvla68Pu93A8y5dfYk3+lGSMMchxwFhN7f32u2eWdwDBHT/4OCXv/3N6OHHPd85+PSjwaVrbtg03zcBMMZJ62oTcm1CyJgQAhkSAReiLEspqz0yABXzvLKjGuElVSIY0aWqJAbYaDvgl1ryXAjTVBFSlEWBRh++poRsOphQLSQg5JxUCXDqqBsn2riUuamRr+YbOSzDZjc7gOpgQgRaK4NEm3+kLwdPc/eaq4jVL2Z2JI3mGA4F8q0rX3/wyQetXt8WFjLUpVJ5yhlmeSqEIIR4tSriuHf91fGTB9n0WRRHK8sSjGtkhKjSfJnaan7EEEutsizJ06QsUlJ5pvVg6+IXt3/VWM5c153HmeX4i9mk3dtCRKU1EY0efjLYv25Li1ly/OizNImBQKxOkjyfPBWUxWWWsDRGXQCgAsIK/dPM9icfvdf75hsiTY7X6/HTB1v7LzDLImW25wFDnC5m0Wx89Rs3bMmB8Zdfef3mj99OOGf5mnRBgAUiIDHz+ZMmonwxHXlhc+/q/NnjUuvp3hWOLccSnmWVmrTST54eeFevSCHSvPjJj37w2h9/x7WkYNBrdd5846/e/rd/XUUnDBCRTPEKWmWz8aeTg2Znq711Sb3w6uj9nzz+4Gc7u1cmT+66luVwzo9GW8O+JQQz1TqA1vrwiweKO1tbO5bgUoDvOq+99i2Wxnc//lVWFJryyaO70egp/8u/fUtp/dHnn9++/dFiepQdPtDZmnN2+evf+vNXrm9327CBbs7bByJKaW0SdETQ2gwim94x6NOGOQCYgrAE0EBgdqjXDPmvkkFMDcKkkBv2jtLKkGq1Ps2vKusnOA1UpBmv9yBvSiXjM6yW+iMNRIxX3EdTRNTyJXU1AQRGr5pxBkBKGQ07rHs+m0oJWZVOmCjChTCpxS+OiqAzXCdrS9rL9Uonq3anzxiURT6eL1q93TKLW0HIpPjs419dfOFl23GTMlvlpT/Y8brbdrvvtAZWdxhneaM77O9c8npbTnvA/HZpu2DZ6Dgo3e2LVx3HO7j3u+7Wbp7ldqOTL6etdo8AkeF0Op5ODveu3LClBMnb3X6utQjb5ATL6cgfXPQ7/ZyJgjEQEi0LpIOWjZZNQoK0dTRpXXxhcfjI7+8li5Nut49MAKAQDIEKVd798OfNnav9btexJENkXnN1/CyOTtzuri5zYEhG74Jx2qxwQdRATtBOZyNKlvM871zYD20nL3IiEEIQUJzlrWbw4e1bv797pzm8cHmrb3GGCJ7v9/avPRsfEwe0HZQWCAmcA+OAjDmOJ3g0PXGGF1ZP7wkplqMD7vmKiJgEIt/zBGemWI/j+IP3fvrqn74Z+rYtOK9oQXxr71I4uPDok4/y5Vyl62Id/T9tJez4PESEmAAAAABJRU5ErkJggg=="}]}
