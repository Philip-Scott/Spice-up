{"current-slide":0, "aspect-ratio":-1, "slides": [{"background-color":"#000000", "background-pattern":"" , "items": [ {"x": -623,"y": 442,"w": 2767,"h": 472,"type":"text","text": "","text-data": "%s","font": "raleway","color": "#ffffff","font-size": 50, "font-style":"regular", "justification": 1 }, {"x": -629,"y": 786,"w": 2784,"h": 315,"type":"text","text": "","text-data": "%s","font": "raleway","color": "#fff394","font-size": 28, "font-style":"regular", "justification": 1 }], "preview":"iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAVmklEQVR4nO3dd3gUVd/G8d9s35AGIQmhGaoIQUCQGppK76DUBykvXRCDFJEiIoj0B5SqAlKioDRBkCTUgJSIlIj0KpLQEpKQZLNl7vcPEAUCHHxUynV/rmv+YTc7M2fOfLMLXGc1EWlgMpnmGo3GfCKiCRHRH+DxeBLcbnc3zWQyndc0LZ/b7X7UB0VEjyGTySQAzmtWq1V3Op0agEd9TET0GNI0TSwWCwzCjx5E9GCa4VEfARE9GRgLIlLCWBCREsaCiJQwFkSkhLEgIiWMBREpYSyISAljQURKGAsiUsJYEJESxoKIlDAWRKSEsSAiJYwFESlhLIhICWNBREoYCyJSwlgQkRLGgoiUMBZEpISxICIljAURKWEsiEgJY0FEShgLIlLCWBCREsaCiJQwFkSkhLEgIiWMBREpYSyISAljQURKGAsiUsJYEJESxoKIlDAWRKSEsSAiJYwFESlhLIhICWNBREoYCyJSwlgQkRLGgoiUMBZEpISxICIljAURKWEsiEgJY0FEShgLIlLCWBCREsaCiJQwFkSkhLEgIiWMBREpYSyISAljQURKGAsiUsJYEJESxoKIlDAWRKSEsSAiJYwFESlhLIhICWNBREqeiljYvLzFy2p+hEegidliFZvNJkbDww6pJhaLVWw2qxgN2j9ydHcymkxis9nEYv53xszm5S12heujGQxitdrEZrWK9u8MhZjMFrHZbGIyGR/wTE18/AOkUKFnxGa5/3MtNi/x9rI9cN+Pft4+JKvVCk3TICJP3FawRHkMHTsN+4+cwsZFE2AxZPc8DUaD4W/ft9nugxr1mmHE2En4dl0U9vz4E+IPHsT2bRsxqGtTGO/zsxYvP9Ru2BKjxk3FmvXRiNu7D/EHDyB2SxT6/6c+tL9wPAGhZTB+/GgE27M7VwMKPVcO3fsOxILIr7Ftxy4cjI/H3rhd+PLzKSiYy+svjIERHd8cgTavVLjncwqFVcLICTMQf+w01s0dBUM2z/EPKogW7bti6szPEb1pK/btP4AD+39C1NpvULdC0b90bcrWboUR/TvBarz7Mc1oRfnwVzBo+Bh8vWotdu75EfHx8di1Yysmj3wDtmzmkGbOge7vTMTpxCQAOr6ZNjDb65s7f3H0fWcMdu0/jP2blyHQmv199UzJFzF83McPmLePz6ZpGqxWK564WATkK4z2PSIQvfMA3B4dbqcDTreOg1HzYb016BqKhFXAoFETEX/yAn7buSTbifqwm8FkQ6WXmmLO4pW4kpoJXdeRlZmK+H1xiImORnTMJlxISoPj193I42O+7WeNZjvC67XCZ19+i+T0LOi6Dkd6Cg7+tAcx0dGI2bgZF1PSkXlqC3wtt9/wfsGheHPoGERGLkb7enffnPlLhiPu2EUAbjQt7Xfrz/OElkTEiPHYe/gMdF2Hrrtx/tRRbNuyCVFR0fjx52PQdR3D2le644ayoFqDNpg7fxE+HvcOcnmZbh8HsxciJkYCuo6tX7x/W9yCChRHpz6DsWnPIei6DpfTAZdbR9yqT25dA7tvIF7t9AbWbt6NLJcHuq7j2pUE7Nm5HdFRUdi0dSccuo4dSz64K5yhpSph7JSZWDR/DioUDbxjLDSEN++FK2kupJ3ahby+N49bMyKsYm2M/2Q+zl5Mhq7rcDszcezQAWzaGIPo6BicOH8Z7rSLqF7c97bX9MpVEJFRe+F2ObBjy2akOYG4b2fBot14PEfOYDTv0APLN2yHw+WB7sqCw6kj4eg2BFtvn7cde72NmF3x8Nwcl7vn7eO5PZGxmL90DS4lpcLtysLRg3swblh/vNSgPa44dcwf1QXe/kHo2Gco1m/7EWkZDrhcTnh0YOfSibe9js0nNzp07Y5n8/kr77t0jebYFPczHE43MlKuYuOapejVsRWeyRsEm9UMTQS5Qsvj2KUMxK36BLabv9X8A/Ohbe9B2L7vCLJcbqRfu4wNKxfj/9o1Q4GQQNgsN6ISXKI6ziRlIjZyPEzajYmfK09BtOs+BAdPJsLlvHEu25ZNvO23WslqzXDw7FUAwLXjm+FtEPjnD8P0hd/iSmo6PG4njsXvwcRRg1CpTAn4envBaNCgGcz4YEEMnGm/oVaJYIgITNYcKBfeAPO+joHD6YbL5YTuSES14kF/jJ1vMMZ+vgYujw7AjYhWFSEGMxq17YulazbiyrU0uJ0OHN6/E6OHvIG6zbsi2enBJwNbwydXCHoPn4oj5xLh0XVcOn8Si+dMRbM64cid0w9mkxEigqptBsGtezCuZ8NbN/szxUpj8JjZSEhKh9PlBAB8+EajP66RwYzmPUbgcloWAGDDvPdgFEHxKs2xZtNupDucyMpIw55t6zGoT2c8WygfvOxWaJrA7BOCTYcScCE+GoG2G6HO4R+IOi26Yuu+k3Bcv4xhPdvioy82wJOVgna1n0f1Bm3x+eLl+PViEtxuF84ei8eMCSNRpfIrOJXmwtZFY2Cz+6Jpu16IXLnh1rw9cmAXxgzth1eavH7bvG3Ysi3y5rkzfo/H9kTG4vTxX7Bk7hQ0qlUJ3rYbN1mzNydD1z34ZuFsHDjxK9weDy6ePYb/jhmC/xvwEZyeLAx4reqtSRdWrRE27T0Kt9OBge3Clffd44N5uHThFGaNH4YyxQvCoN3xHM2MUfM2AHoWejauhNqNXsOshd/gzIXL0HUdVxNPY9qYwQgrmv/ujxkGKyYtjYXbmYpOdSugTrN2+DRyFc4l3ohAwpl9GD9tAdy6G8Nfr3XjAhrNqNf+LVy4lg6n0wnoHswY0h4FSlZFVNwpeFwObN+wAq3qhcPXy3LX+RQLb4NUp46tX01GqecrYMCIj7Br/+EbkchKw5JZHyHudApO7V6JXDdvoIACJbFs0164XC64PTqSTuxAoTxB6DVyJtKzdCQnnsMXM8ejXvUKyGG98Vu9w7tzoLsc+HLBHPxyJgEejwdnD+/D2z3aI1/g3bG25XwGsUcv4drZH/FiqefQvtubWB0Vi6TUDOgeN36KXYkFq7bBk56ImsVv3Fwmmw8ixn2O61lOOF1uwJOJNtWKoGrjLjhxIQ2OjBR8OXcSqpcvCYvxzo9pGjq8MxNujwuT3mqLCuF1MWHGfBw5fR5uj46MtPPo3LAiStbqgGsON5IvnMCe/UfgcHngSEvGhq/n4bWGtZDLxw4RQZkmfeD26Ihe8QW27T0MlwdIufQbIudOQYMaL96at68N/PiPeXv8V7hcTlQPr/bI77GnJhZ+Oax33GR2LNpyGACg6zoObl+P7u2bI8jXBhHB4E/WIOPqKZQKtMDunxejpi/GtUwnUhJPoHebOjAb1M/bZLHD3yfHPR/3yheGo1eyAI8DSSnXoQNIunAKiz/9L9q0aIzQ4Hu/i/EpVAnnrrngcWciOTUduq7j8q/HsWDWJLzWrBFC8+bFwo0/I+1sHIJtGmy+wRg9cykyXB4c/mEtZi+NgsdxHV98NhcJyelITzqHfu1euc/fm2gYPm8jACAlJRkujw5PVjq2R63CgN6dUa1CaVRo0hduXcd7nWpDxIDK9Tvg0K9X4Ei7jInvj8ZFh44DW9dg3faD8OhuxHw1HaHBPndcnxxY+ePZW9dn7+bV6NK6MXJ7W+85FuVavQ0PgMz0VGQ4nNA9bpw4uAsT3x+Mhq/URL7Q53H4Uga2fzUJFoMguEg5LNu4F7ruxup507Dp4BlkJhzGnEWrcd3pxq+HYvFy+SL33J/B4oOo4+mA7kLytRTouo705ItYGfkpurRrhbCi+SEieLnbB7c+yu3dth6D3uiKF54LveP1DBg1Pxq/O/dLHCK6/weF89xx7Q1eWPrDidvmbacWdWC3GB/5PZbd9kTG4q4L7V0AOw5dwC+7Y9C+YTjMf/6tYfRDzLHLOLF9OTr2HoKj56/ClZWO7xZ/jKJ5/P7+Y7H54/3pC/H92pX4YNjbqF2lLOwWk9LPGr1yY/zsL7Hu2+UYNTQCNV4Mg838x88WfKExrma6sWTSILTs1A8/nbgAV9Z1fPnxSOSym/DmhKXQAXhcDmxbG4nKJfI/cJ9Vm3RDVHQ0PpsxGR1bN0HeAF8Yfp8HRjtmrd2LtPP7Ue+lOvh40Vpkujw4E78D9SsWR67QKkhId0LXdSSe+QUj+rSF1Xj3HDL6FcX+U5ewP3YdWtetDJNCnANCy2Pp6u+xPHIB3urdGaWLFoDxT9e18RsToOsuDOhQH/1GTMZvydeRnpyAET1bwmrLieU7jgIAMlIuY8mMMcif696BFxGIZkKPYdMQtX4tpnw4Ek3qVoeP3XLXuz+z3Q9NX22DF0o8A8O9zsNkx5KYozhzaDf6dWwKb2v219/oE4q4o4nZz9vHcHsqYiEi8A8IhLft7rfZ5sByuJDsuPGW2ZWF/du/x6uvVMzmbejjv1VuMRBuXcf1tDS4XU4c2r0Rbf5081m9c6JS1XCUKl4IFtP/fn6GHHmwOf4yXFkOpGc6kXL5N8z9aAjy+N/8VxPNgEIlyqBqpfLI7e9939fKlTsIXlbz/3xMv2+D/rsWgAepqdeRlZGGjSsWoNJzBW89njO4IKpXD0do3qC7Pyr+C5u3fwD8vG0PfF7O3EHZztvHcfs9FprVaoXT6RQA8lQx2qXbWwOleIBJYjdukI2xuyXD6XnUR/WX2PzySI8+vaWAn0F+2BwtMdt2Slqm6x/co0Eq13tVWtevIuePH5R169bLkTOJ/+D+1OUp+oL06dZetPRLErX+O9m17xdxeZ6yufuY0TRNLBaLPL2xIKK/xe+xeCr+BycR/fMYCyJSwlgQkRLGgoiUMBZEpISxICIljAURKWEsiEgJY0FEShgLIlLCWBCREsaCiJQwFo8bTZPgYB8xPeSVsVjNYry1IrYmuQN9xGq6fYlszWiUoCBfCQ7wkn9pIfFbrHar5A3xE78cf201a5PZJJY7zkc0TXIF+EhIsPc9x8tsNT/0WFL2OIwKNKNJylcpLtXLBt/6s/wlisjXS7pIXpuIwWSSos8VlP79XpZCAaZbz/EL8JWGLSpJ58ZFlfbjFxwos+b3krjYofKf8GDxy+0vjRqWlmCfm69pMEqniJbyftfnRUTEbLVImQrFZOz49rI/bqi0qBokNl9fGT35ddkT+46893opseWwS+165WTGzM6yPeotWRXZXTZFD5Thr5e4cW4Go4S9UEReqpjv1nEEhRaQZd/0liLe9y+K3ddb6tQLk9Cgm8veawZp1LGuzB1e88br5AuUzj3qyPKv35At3/WVb5b0kLgt/aVsfquIiNi8c8jLdUpJ0RCvmz+vSc3mNWTh2Do3TvfmuA58t4Xs2TlM3nn9OTFZLVK+SgmZMLmDbI2KkLVLe8j6NRHy+Xvh8vvRmixmKV2+qIwe107273lXXquRR2n86f4YiwfSpOfgV2XZZ6/LlIFVRRORsCrPy3crusuz3k4JqlBatmwaIF/OaStD+1YViw6x+XjL+590ki2re8uUMc2kYnE/0TRNyoY/L6P7VpXsbkHvwECJjOws106eF0dmuoRUKCsx6/vJ/Dmd5KXnfMRst8vAD9rL7JE15eKl6zJgTDvZHh0hU4fWkHM/n5aUTEjOAnll9cq+EpiVLMkZWeLxzyObNkfIwA6lJHbtLmnTbrbUbDJbDiU6JDlVl8YtK8uK5X1lxaLOMndkLdFEpFi5ErJ6RU+pHqKLpXARGdyzgmT7LRnmHBK5rLcsnN1JWlfLIwajSbq+3UKWTGko166mSs9BLWXzyq5SPp9Rpn60Suo3mS4dBn0vmZlZYvbPLf0iGssPG/vLormdpOPLBUQzGqV1j4byzewWknY1RVr1aiCx0RHyxeTGYriaIKeTPGK0+sjSb9+Uae/WlGO74qVLl8+kVsPp8t2+a5J0NVNq1Ckrc+d3kx3RA2T6sFqScOSMJGfq4hcYJAO6Vxb7g74ahO7LaDKZRnk8T+aiMP+WhHMXJX/ZZyVmWawUe6mqTImoIOcuO8Xfxy7N6xaWiaO+ls+jL8uLwU7ZnmiRhZ92EMeRY9J38Gop/VIZWbN4h7Tu11wGty0mCxbskBMJ6dnu59Cuw5LsXVA61CkgKVeSZcHyo1K+kEFmrj4vk6Z3lFA9TfIWyyVBhQuJb+oFGTJspUyY/YNcEl8Z2r+GFAuyyadTv5Pvj2vSv0MpcWZkyCdTv5NRk2Ml/vgVSU13SUipYvLhgHApXDhIvA1OWfvtT5LqFSB71u2WwPLlZMaw6nIuMV18vazSomlJWR25Uw6dS7v7YHWPHDp+TWpVCpSZi+NlyLiOUjNYF68Qf/ENCpZnfTKkY5cFsnjtUTmXkCZZLl3a9KovLaoWkLCwEEk4eV4iV/8iYWFBMmv+XnlrdAdpWsIq4uctPoGBUjEEMnzkahk9ebPsOpIpY8c0klIFfGXFF5ul/9C1sufQRUlOzRKLXy6ZOqmZhIbklHy5jLIl5pDM+2yTfDRzh/zmzCHDBtSU4iFesjH6Z9l/PEm4asvD0zRNjEbjk/0lQ//aZvbBviMf4uddQzB/QkOE+JlRtHRhdHz1eeS++f0gzfq2xOWToxHzVSdUDwuAJgKbf04cPDURB2MHYlSfivCzP3hBVoPRALvVBE0E9To1wKVj72NXdF90algEJpMZLdpWRs0X8sD4pyXjfINyo36NUFhuroOpGTTYbSZo2S0rp2nwslv+WH7PZMf3P7yHw3veQeS0pgjNbUWBZwuiS7vyCPG//7JvYbVeROLJMYjbHIGI9qVgNhpRr2kFNKoRCnN2a3KajPCym2G8+T0ZxSqWQcKpsfhx6wAM7lQGdrMRNeuXQ7OXC986FxGBweqFZg1KwNua/fjZ7BZYzXc/5pM7AA1qFbrttbg9/Pb0L6v3NwvOm1OMbqckXEqX7EbK5m2XYH+LJCSkivP3Zd40TfLmyymO1OuSlOp86H2abVbJH5xDrlxKkbTMf+7dX0Cwv9g1t1y4eF30h5gGBrNJCoT4SkpSmly7/vDL/BlMJsmf11euJ1+XpLSHHx/6d3BZPSJSwmX1iOihMBZEpISxICIljAURKWEsiEgJY0FEShgLIlLCWBCREsaCiJQwFkSkhLEgIiWMBREpYSyISAljQURKGAsiUsJYEJESxoKIlDAWRKSEsSAiJYwFESlhLIhICWNBREoYCyJSwlgQkRLGgoiUMBZEpISxICIljAURKWEsiEgJY0FEShgLIlLCWBCREsaCiJQwFkSkhLEgIiWMBREpYSyISAljQURKGAsiUsJYEJESxoKIlDAWRKSEsSAiJYwFESlhLIhICWNBREoYCyJSwlgQkRLGgoiUGEQEj/ogiOixBxOARJPJFOJ2ux/1wRDRY8hkMonH40nQRKSByWSaazQa84mI9qgPjIgeK/B4PAlut7vb/wMRdrD+bfFS2wAAAABJRU5ErkJggg=="}]}
