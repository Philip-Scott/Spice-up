{"current-slide":0, "aspect-ratio":2, "slides": [{"background-color":"#ffffff", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/beige-paper.png" , "items": [ {"x": -522,"y": 442,"w": 1410,"h": 509,"type":"text","text": "","text-data": "{title}","font": "raleway","color": "#000000","font-size": 37, "font-style":"regular", "justification": 2 }, {"x": -560,"y": 906,"w": 1447,"h": 315,"type":"text","text": "","text-data": "{subtitle}=","font": "raleway","color": "#505050","font-size": 21, "font-style":"regular", "justification": 2 }, {"x": 1096,"y": 374,"w": 715,"h": 816,"type":"image", "image":"jpg", "image-data":"/9j/4AAQSkZJRgABAQEASABIAAD/4gxYSUNDX1BST0ZJTEUAAQEAAAxITGlubwIQAABtbnRyUkdCIFhZWiAHzgACAAkABgAxAABhY3NwTVNGVAAAAABJRUMgc1JHQgAAAAAAAAAAAAAAAAAA9tYAAQAAAADTLUhQICAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABFjcHJ0AAABUAAAADNkZXNjAAABhAAAAGx3dHB0AAAB8AAAABRia3B0AAACBAAAABRyWFlaAAACGAAAABRnWFlaAAACLAAAABRiWFlaAAACQAAAABRkbW5kAAACVAAAAHBkbWRkAAACxAAAAIh2dWVkAAADTAAAAIZ2aWV3AAAD1AAAACRsdW1pAAAD+AAAABRtZWFzAAAEDAAAACR0ZWNoAAAEMAAAAAxyVFJDAAAEPAAACAxnVFJDAAAEPAAACAxiVFJDAAAEPAAACAx0ZXh0AAAAAENvcHlyaWdodCAoYykgMTk5OCBIZXdsZXR0LVBhY2thcmQgQ29tcGFueQAAZGVzYwAAAAAAAAASc1JHQiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAABJzUkdCIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAWFlaIAAAAAAAAPNRAAEAAAABFsxYWVogAAAAAAAAAAAAAAAAAAAAAFhZWiAAAAAAAABvogAAOPUAAAOQWFlaIAAAAAAAAGKZAAC3hQAAGNpYWVogAAAAAAAAJKAAAA+EAAC2z2Rlc2MAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAFklFQyBodHRwOi8vd3d3LmllYy5jaAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABkZXNjAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAC5JRUMgNjE5NjYtMi4xIERlZmF1bHQgUkdCIGNvbG91ciBzcGFjZSAtIHNSR0IAAAAAAAAAAAAAAAAAAAAAAAAAAAAAZGVzYwAAAAAAAAAsUmVmZXJlbmNlIFZpZXdpbmcgQ29uZGl0aW9uIGluIElFQzYxOTY2LTIuMQAAAAAAAAAAAAAALFJlZmVyZW5jZSBWaWV3aW5nIENvbmRpdGlvbiBpbiBJRUM2MTk2Ni0yLjEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAHZpZXcAAAAAABOk/gAUXy4AEM8UAAPtzAAEEwsAA1yeAAAAAVhZWiAAAAAAAEwJVgBQAAAAVx/nbWVhcwAAAAAAAAABAAAAAAAAAAAAAAAAAAAAAAAAAo8AAAACc2lnIAAAAABDUlQgY3VydgAAAAAAAAQAAAAABQAKAA8AFAAZAB4AIwAoAC0AMgA3ADsAQABFAEoATwBUAFkAXgBjAGgAbQByAHcAfACBAIYAiwCQAJUAmgCfAKQAqQCuALIAtwC8AMEAxgDLANAA1QDbAOAA5QDrAPAA9gD7AQEBBwENARMBGQEfASUBKwEyATgBPgFFAUwBUgFZAWABZwFuAXUBfAGDAYsBkgGaAaEBqQGxAbkBwQHJAdEB2QHhAekB8gH6AgMCDAIUAh0CJgIvAjgCQQJLAlQCXQJnAnECegKEAo4CmAKiAqwCtgLBAssC1QLgAusC9QMAAwsDFgMhAy0DOANDA08DWgNmA3IDfgOKA5YDogOuA7oDxwPTA+AD7AP5BAYEEwQgBC0EOwRIBFUEYwRxBH4EjASaBKgEtgTEBNME4QTwBP4FDQUcBSsFOgVJBVgFZwV3BYYFlgWmBbUFxQXVBeUF9gYGBhYGJwY3BkgGWQZqBnsGjAadBq8GwAbRBuMG9QcHBxkHKwc9B08HYQd0B4YHmQesB78H0gflB/gICwgfCDIIRghaCG4IggiWCKoIvgjSCOcI+wkQCSUJOglPCWQJeQmPCaQJugnPCeUJ+woRCicKPQpUCmoKgQqYCq4KxQrcCvMLCwsiCzkLUQtpC4ALmAuwC8gL4Qv5DBIMKgxDDFwMdQyODKcMwAzZDPMNDQ0mDUANWg10DY4NqQ3DDd4N+A4TDi4OSQ5kDn8Omw62DtIO7g8JDyUPQQ9eD3oPlg+zD88P7BAJECYQQxBhEH4QmxC5ENcQ9RETETERTxFtEYwRqhHJEegSBxImEkUSZBKEEqMSwxLjEwMTIxNDE2MTgxOkE8UT5RQGFCcUSRRqFIsUrRTOFPAVEhU0FVYVeBWbFb0V4BYDFiYWSRZsFo8WshbWFvoXHRdBF2UXiReuF9IX9xgbGEAYZRiKGK8Y1Rj6GSAZRRlrGZEZtxndGgQaKhpRGncanhrFGuwbFBs7G2MbihuyG9ocAhwqHFIcexyjHMwc9R0eHUcdcB2ZHcMd7B4WHkAeah6UHr4e6R8THz4faR+UH78f6iAVIEEgbCCYIMQg8CEcIUghdSGhIc4h+yInIlUigiKvIt0jCiM4I2YjlCPCI/AkHyRNJHwkqyTaJQklOCVoJZclxyX3JicmVyaHJrcm6CcYJ0kneierJ9woDSg/KHEooijUKQYpOClrKZ0p0CoCKjUqaCqbKs8rAis2K2krnSvRLAUsOSxuLKIs1y0MLUEtdi2rLeEuFi5MLoIuty7uLyQvWi+RL8cv/jA1MGwwpDDbMRIxSjGCMbox8jIqMmMymzLUMw0zRjN/M7gz8TQrNGU0njTYNRM1TTWHNcI1/TY3NnI2rjbpNyQ3YDecN9c4FDhQOIw4yDkFOUI5fzm8Ofk6Njp0OrI67zstO2s7qjvoPCc8ZTykPOM9Ij1hPaE94D4gPmA+oD7gPyE/YT+iP+JAI0BkQKZA50EpQWpBrEHuQjBCckK1QvdDOkN9Q8BEA0RHRIpEzkUSRVVFmkXeRiJGZ0arRvBHNUd7R8BIBUhLSJFI10kdSWNJqUnwSjdKfUrESwxLU0uaS+JMKkxyTLpNAk1KTZNN3E4lTm5Ot08AT0lPk0/dUCdQcVC7UQZRUFGbUeZSMVJ8UsdTE1NfU6pT9lRCVI9U21UoVXVVwlYPVlxWqVb3V0RXklfgWC9YfVjLWRpZaVm4WgdaVlqmWvVbRVuVW+VcNVyGXNZdJ114XcleGl5sXr1fD19hX7NgBWBXYKpg/GFPYaJh9WJJYpxi8GNDY5dj62RAZJRk6WU9ZZJl52Y9ZpJm6Gc9Z5Nn6Wg/aJZo7GlDaZpp8WpIap9q92tPa6dr/2xXbK9tCG1gbbluEm5rbsRvHm94b9FwK3CGcOBxOnGVcfByS3KmcwFzXXO4dBR0cHTMdSh1hXXhdj52m3b4d1Z3s3gReG54zHkqeYl553pGeqV7BHtje8J8IXyBfOF9QX2hfgF+Yn7CfyN/hH/lgEeAqIEKgWuBzYIwgpKC9INXg7qEHYSAhOOFR4Wrhg6GcobXhzuHn4gEiGmIzokziZmJ/opkisqLMIuWi/yMY4zKjTGNmI3/jmaOzo82j56QBpBukNaRP5GokhGSepLjk02TtpQglIqU9JVflcmWNJaflwqXdZfgmEyYuJkkmZCZ/JpomtWbQpuvnByciZz3nWSd0p5Anq6fHZ+Ln/qgaaDYoUehtqImopajBqN2o+akVqTHpTilqaYapoum/adup+CoUqjEqTepqaocqo+rAqt1q+msXKzQrUStuK4trqGvFq+LsACwdbDqsWCx1rJLssKzOLOutCW0nLUTtYq2AbZ5tvC3aLfguFm40blKucK6O7q1uy67p7whvJu9Fb2Pvgq+hL7/v3q/9cBwwOzBZ8Hjwl/C28NYw9TEUcTOxUvFyMZGxsPHQce/yD3IvMk6ybnKOMq3yzbLtsw1zLXNNc21zjbOts83z7jQOdC60TzRvtI/0sHTRNPG1EnUy9VO1dHWVdbY11zX4Nhk2OjZbNnx2nba+9uA3AXcit0Q3ZbeHN6i3ynfr+A24L3hROHM4lPi2+Nj4+vkc+T85YTmDeaW5x/nqegy6LzpRunQ6lvq5etw6/vshu0R7ZzuKO6070DvzPBY8OXxcvH/8ozzGfOn9DT0wvVQ9d72bfb794r4Gfio+Tj5x/pX+uf7d/wH/Jj9Kf26/kv+3P9t////2wBDAAMCAgMCAgMDAwMEAwMEBQgFBQQEBQoHBwYIDAoMDAsKCwsNDhIQDQ4RDgsLEBYQERMUFRUVDA8XGBYUGBIUFRT/2wBDAQMEBAUEBQkFBQkUDQsNFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBQUFBT/wgARCAMOAjoDAREAAhEBAxEB/8QAHAABAQACAwEBAAAAAAAAAAAAAAEFBgIEBwMI/8QAGQEBAQADAQAAAAAAAAAAAAAAAAECAwQF/9oADAMBAAIQAxAAAAH3cpQCgAEAAAABACgEABQAAQAgBAQHE+Z84+9cjkAAAADkAAAADLmIAKAAAAAAUgBCgAEABQACAEIUgIQhxPnHyl+1n1rkACgApClIUAAAy5iCgAAAAAAAAAAAAgBQAQAHEAFBxPnHzX4x2LPtQAFABQACAoKCAzBiCkKAAAAAAAAAAAAAACAAhAClKQ+R8peafWuZDiCAoBSggICgAEMyYkAAAAAAgBQACAAAoAIAQpCAAoKCAHIpDgQgBSlKQEAKUhSAzBiQAAAAQAAAoAICAhSlAIACEAKUgKAUAA+ZxIReaUFAABQAAQzJiCgAAgKQAhSFBQQEIAUpQCAA4gApSAFBQAQ4nzIQ+hQUAAAAAAzJiCgAAgAABAUAAEIUFBQAQAhClKCAAFABxIUhCkBQQoABSAAzJiCgAEAAABAUAgIClKACAAA4lKUAEABQCA4nIoIcSkIACgAAAzJiAUgABAUhQAAADiAUoAAAAIUFABAAAAQhSgpxKQ4gAoAAAMyYgAEKAAQoAAAAIQpQAACAoABQCAAAAEICgoAIQAAAAAzJhwACgAAAAAAAApCApAUAAAAAEAAKCEAAKUhQDiAAAADMGJIQFBQAAACApQcSlBCEKCHIgAKACAgKQoABAAClAAIQAAAgMyYcAhQCgAoBAClIACkICkBSAAAAgAAKAQAAApSFBACAAgAMyYcgAKAAClBAUFIAACFAABACAAAAAFAIAAClBAQFBAQAAzJhyEIClBQCggBSlIQoABQAQAEIAAAAAUEAABSgHEAApAQAAzJhTiQhY5VyKAAAUoBSAAAFABAADiAAAACggAABSkBAAAACAAzJgz4S8inNPpXIgABQCgAEAKACgEABCAAAAAoIAAACkABCgAAEAMyYGOVcgU5gEIAUoAAAAABClICFB1zVTUTCy44+h3k2CtxNlOQBAAAAACAAoAABAZkwkc6hTkUEBAAUEKQpCgAAAAhDWo8eXCY3OS7LLt0cS11TTzEWaplN7uPrhmKAAAAAgICgAoAIDMmKIQHIAgAIAQoKAAACAoIY88FlxmGXoON3mzQMcvkfHDPBHKtgjG5Y7LZtOWPn66JnjvVx9prmCFAABACAAoKQAGZMWQEBQCAEIACgAFABAAatH5vmXsmGX2Ohrz85lwOePxyx6OWPwsp2McvvLkcctlwy3PPDOZTTK1bPD9IpkaoABSAEAICgAAGZMUAAAQAEBAACkBQUEIU1OPzXMv0Lry1ldQ156Jt14nZrAAHGucQq7Dp2bTMvQssMVXnWzD9P2d4AApAAAQhQAAQzJigUFICAgKQEAAAKAAQx8fk+Ze+a89dTz7HPSd+ngnKXjXGywAoWWnBO3jlsuGfrlmsmC2a/0xVAAAAAAIACAGZMSClABAAAQhSAAHIEBAfnOXNYZZvHLyvDLSujRVscaliAAAKvKXhcfvLverb6dZ5Hnh7Rlj6LQAAAAAAEAOIM0YgFKUEBAUAhCkAAKUgIYA/M2OXt2vPzLHLz3dp4LxOGWKAAAAFI+ky42dvDL2PHL62edbNf6woCwoAAAAAQEBmTEAFAKAQgAAAAAAAPEIwuvZs8eO5TFV8MsYlWIBVECKQAOcyptmvL2qvB88P01ZslAUAAAAAEBCGaMQAAAUpCAAAAAAAA/LMega9mOxvjuzDgcMpxQDlMhLB9Mcuzhs6mzVxsiKFl5S5PG+zS6hljvmePq4BQAAAAQAEIZoxAAAAKUhAAAAAAAD8hy+3atnl9aNZ1s8BEq/bHP4ZYLAMnp3ZPVnrPXzWUSxCuUuQxy9Vxy6FxzGzD3CLQAgi1AAAAQAzRhwAAAUAgAICgEAAB+RJfYtWzzOzTK+GeEKc5dk4+3V+7gEBsfL0d6XT+vmFlgsRV+8y9UwvRszuzD3YAAAkKAAAEAM0YcAAAAFIACAAACAofk6PQdW3UTRcsfhnjEq2PSPN9Dzj0vP4ZSA27k6frcdN6tAHPHPhcSDtTL1PHLA3H0TPH16FBCoWJSFAAQEKDMmIAAAAAAAAJCkKAAH56jpa9nHHLzvPD4Z4xKpPVvN7/ADfv5Ohs1wG8cnR8csdN6dNOzr2drXvxm/kAyOOfrkvmeWH6Ts2woqCFAACAAAAzJiAAAQAoAAAAAIAAaLHgGOW669nm2eONzwollnq/n9mi9WjA79Ih6BxdOP269Q6NQ2Xi7ensww3RyirtOvP0A832a/12c6QFAAAQAAAEM0YgAgAAABQACgpDjAtAQ/KEblp26bbqGzVxonYw2ek8m7XdmOodfOB6Nw9WE3atU6NQ9K8j1dB9Pz+nnrJ3Jl6Dry17PH1zLH1igAAABAQFAABmjDgEBCgAhSgAAoiUAAhWnx+cZd41bfOc8cXngNm4u3YstXxl887eUI9N4erW+jVq2/VY9j8T2PG/b8glXcNeeXsxeeH6pORRQAARKAAgKAUzJhwQAAAAFAIUAAAoIAePx5XhnmtezRturpZT0Tz+7rb9Gc0bPJ/R4wX1Pz+vVOnRq+7XmNG7fvP7fKfX8sZvDPaMWubcf1OmYBRQCBBQAEKAAUzJhikAAAAAAALEFUAQFADxmPJMctg17NU2a914unobcNy593inpcXFC+r+d2ar06dT6NO8ef3fa46F38WwYZ5MxmeH6fM8UAChIACgAIUFAMyYYAAAAAAQoAACgAQFIHnp+f1+2vPbubf103TRs8B9TihT1Pze7Xd+nTuvn9d8n0tQ7OXrbtXwyx2/LH9BneLQAAghQEKAAAWFDMmGAAAAAAAAAAKASFAIA6Z5CaHq2bjx9Ww6Nng3refjMpT1/wAztx2TSO3m9m8f0fFfZ83bs9fsxu4KBSFIEBKoAAi0EKEKZgw4ICkKAAAACFgBQsKgBItABHCPNPO7u3qz8N9Xg1TKVfY/L7e/o6NL7Ob0rk6fQva8jKAFFICkKRBQAgKCggKQGZMOQAFhQAAAgABYUBYlBAUAEQ0HzO/7a74j6XJo+3WX23y+zYOXp+cyzvXz7z6nnSLShCwAAOIqgAEKUkKAQMzWGABQAAIUBAQFEWgEWhAAAAar5/X0OXd4V6fJp27VZfdPO69l5t9jO9/Ns3byCwyFSKRIUBKohQCFCkBCkKZkwwAKAAAAQAEEWhQBACgAAMNx78JxdPgXoc2odGjlMvevO69n59qXZfU4svu0y2pQsS1BAUEKAQoIVSCFCFMyYUFAKCAFAIQoBAWLQAAAAAHQ59muef1+Rd2ny7p5+Uv6D83r2DRtku4exwdvPCRbKKRACUKIlUAAoECCgBmjCghQABCqAACEBRFoAAAAADq6c9b8/s8i7efyro0/THL9XeZ14TR0d247r7Xm/W4gCgAlIpKQLSALQARKAAzJhgAACFAKIUAIIFFBAUAgAKR1teWB8/r8A7NWj9Gj645/qjyuzq6tnGt49rzOdgUikFBFJVAALCgAESgAMyYYAAAAhRFFAABCkKARAACgHV1Z6553X+fe3Tp3To7GOf6n8rs6evP6G5ez531yxi1IFFRVhQACLSFAACAAGZjDUAAIUEByAAgBQAAARAAUgOpp2a7wdX5y7dOtdHP2cc/1d5nXitG75LvHs+b2M8QpICglKSrCocgCQKKEBACRmjD0AAAABQCFhQCFICkKARAAQx/PuxXHv/M/bp17fp7uGf6q8zrwend2k3H2fO++eJAW2IgUEpSVRAUAIUAgiUjNVhwQoAAAhSFBFIWgAhQCUipAVIGL5d2M5t/5l7dGE3a+7hl+qfM6sdq2ytu9bz+1swChYEFAWFBCgAIUCAqRBWaMOCFKCAAQFQogKRaCFABChxECCXF8u7Dcu/8AM3oc2I26u7hs/VXmdfQ07PrlNl9bg7mzBVIXEpUKQAAoIIEBaQoSFDNGHBClAABAAIAUEKRQABUBIggYzl367y9H5/8AS5NW2a+1hs/V3l9WM07u1cdi9Xh727WoIoCxKSggKQIAKAACVYjNGHoAAAUgEWoItSAFIlWBSFICEhbZIuJ5N+r8vT+fPU4cHnh9sM/1b5fXi9HR92Ozetw5HfqAqCwoQoIWpEFFIgKFIIAGaMPQkWgAAIAUCAoABFBACEVFspDD8XToXPv/ADv6vBZfpMv1D5XXdW2VsfpcWT6dIBOQAAIKpIgpCkBQSrAlWIzRh6AAAAgBQABCkBSEKCJQhQWoa95vX5ncvD/Q4+KfXHP9Oed1dzn3cJc76HHl+zQEWy0JCkUi1IAKgAi0hbEAAzRhyEBYtAAAAAQAoEACABSAU4mueZ2aDunhnby9Y+mOX6N4OnP8+3545ZTr58738gUqiLSFCQAKKEiVQAQCFIzRhqgUgoABBCrFoCAogCUEARQKlr4a8tf8/r1Dow/P/XzfIuOXvXD0bbzb/nryynXo2H0eJQKTkKRKQIpKWhCkBAAAIi5tMLQAAAAQBRQohQhREFSUAIAtnT0bNT4evyzr1eX9PPxs+ky9i4On0Dk36Vuw37G7b6/nFIKC0iAAFoCAkAAAKkFzcmFyAIUgKARCikKpCgpAIikAAKipiuXfoPD2+F+v52KyiOS+q8u31nj6PE+7n9f8zt3f2/LtlAKKghSBahQSIBSABFIVGbswgUiqCQtSKQKAKCFUQBAAqwJSBLrPn9flE2ePen5/KXjZ9sM/SNOftXD0aN145fg6d99bze3sxqWpCrEpAAUAiUgKkBagQsSs5JhFUCWpKAEi0VAAoIoIqwIKAABxxa35/Xhtjr9vJ+aqlc8ct61Ze8ed1Yjpx6PF07/6nnd/fqUJAFIKKkUgKCBAohUEAM2YVQCWpAKAAssAKSkpBQQAUhSFHU1Z4Hh6eHTq1Do0+GV1LGOWzYv0f53X8OjDVfP7/QvS8zK9eiEAAAFIAEAUAQAkCgzZhahYUS0gQKAKgUKBEFIKsCCkBSY/m3apx9Wz+hx+f54/nuz5Wc5nlo/UHmdfxzmt8fdunf52c9DlRxUgAhQCSrAVAEpAgAAM2YawRaEtAIgKSrC0JLSFQQCkUVIUAmF4ujVNHR6F6fB41MvF7OrZZl9E/V3l9mqsu5y79h6+bZfV4UQAkKAKRKoJIoEABCggM4mFtqRaAlFIUlWBKpBAAIoqAABSIuueb14rK7x38ficvk9Yi485nwuP6q8rtw+3HyHonu/Fs3H1eEgChIpBKBKpBEABCgEAM4mFtCKKIKLSUEAVJFQoIEqpQSrAgl+ON1/g6urtm4dnL4rL4hlJLzl+WWP6Q8jv2jbhgNz78O/evZ8znYAApElgCARRCgAAEAM5ZhFoALCygKsCApEVEAFllACwJSF6GnZrvJ0d7o1bF06PzzLpS4HLDnjn8ssffPM7d4Oxvw17zezd/Z8ztbMFlABBHG2xAQApQhQIUhAZxMLaBItIosooBCkQKiFIBVhSAABhOXfqnJ07z6XF3M8PB5l47ljD645fLLH9CcHVuuvLu9unzzwvY9C9nyMv06FgKQogiEAABQUAAEBm0wigUCiF5JApBQRQiFAoIAIUCGucXTqmnf6b6fn8D83S4BdZyx545cMsfbOLo9I59uwelyedeD7O5er5eZ6+ei0QFJEAAIUAAoQoA4mcTB22ALSFEqpAtCFBCgCAFgihAX5y615/V0c7u3dx8T89y+VZQfSZcLj6xy7/AFvi35/0uPRPF9bZ/Q4M53c1SW0hSRCkLSCRQAAKQAEM4mDUUopIUBYlIFoQBSFsKgSiJagi9PVnhePo6u2bh2cvSPzOuMxuuZ4/THLhlj69z7fV+Ho67LHcvRmevl2X1OIAKCBC1QREsABCggABnEwS0pyRbECUBSJVgAgKS2hCoAAIx2jZr3L0Zfq05zfp6R+epl5rljTnMuFx9y59vovF0eW7Lm+fbtSbf7HmgCghQKsktQIACAAhQDOJg1oKC1EKiAApAUItRQiixKCSwGG49+taN+8ejx9jLHAn51mXzjT88fpMuNnrWrP17g6On06vE9z0/wA7q9E9Pg+uWIFAAAAIACAEKAAZxMJaECirJLZAEKAUItFEgUlWFkCA1nzuvE3LffQ4qYQ8Al8+yllpxs9W17PXvN6u906cPnli/N6919Xzu7u1gCgoBAAQAgAAKAZyzDLCQKikS1AAAFBCirEFIWIigfDDLXfP6untm7d3INaX84kjWsnKXim94Ze4+b15Lfq+2/DVPI9DavU4Mn1aAKACgEAIACApQADOWYWCwAAgABQEKAKEWogBADG6NuK5d3z3Y7X18w19fzsa2dWrLwuPpWvZ6h5nXntuvNd/Nofg+ttXp8GY7eYCgAAAgAAAKAQAzhhiAgAIAUAAAAoAIQAAwvJvwujdnuznyu7UNcl/M1dQ6y/NIegYZeh8HVtWLaPU4tC8D2Nh7uLO+jyAUgAAAAABQQAAhnTCkBCkAAAABQQAFICApAa9wdWD1bd59Ph+lg1c/Ny97HLXa+mN+lm8Y3eubdumu570OXz/AMT1u/lr3P2vMpAAQoIUAhQCkABAUzhhAQAAAAEKAUhAACAFBxl1DzO3G5X0T0uD4y8q13DL8/69mRxZbHLnMvphkzx3fTlsTHv9ejXPP7vli3j2fOIABAACkKAAACAAzpgwQFAAIACggAABAUFB19eWG5OjqW7F182O1bMLjnrOrZ0ccuUvIyjHZJjkcscZhs7zHG69n2KbJ6vD2c8YAQFIUAEKACAAAGdTBKAKCAAhQUgBAAQFKClMXzbsZzbuzsxwUy1vXszLHNJyyxwec1/Oa7k1/Jgcp6Dpy9i5c/J9zN68tu589j9Ti72/UAIClAIQAAAAAEM8mAWgFIAUAoIUAhAQFKAciGE4ujoaNvx3Ya9WvZNfzmu544fLHZI1jLH4ZYw+sz3rTn7rw7vM7u8u6tfpemewbdGU69AoABQCEAAAAAIDPWYCUAADkUAAApCAgBSgAhrPmdvm+/Dybfj188PnceNx42EycyxlxL9JlDZ9d/RXndXnW2+PdWr1jze71Xq4c33c1AKAACAhQAAAQAztmAlAFBSlAIUAoAIACkAPhhlrPm9mi5bMFnPMu7jlkT53GZYwAsVc/o3fpXg3aLvw8L7Nftvh+r6B18OxenxgUoABCAAoAAIAQz1mBlEBSlBSAAoAKUAAgBDH6NuE4enxy9Ot7ccL1cXX2auNx42SznHChDLYZZTR0/ozjy1vZPBO3V7f43o7Vt59n9fgoKAAQAoKAQFIQEKZ2zBywhQUpACAAoKClIAADiYfi6MFo3+IdE1Tq5vncJUTjZLAALLyl/U3mdfzPPfQ5988ru7GM2v2PP8ArlKUAEIAUAAAAEAM8mCUQApQAQgIUFBSFAKCHE1zzezAYbds9Di0LJ46uByw4Z4xABQQsv6W83rzeGXZ9Lk6XndnT59u0etwd7brFABCAEBQAUAEAM8mBUAClIACEABQACgFIfOXVfK7sNcvQ/V8/knwXzHHLx1lgs9fG4iyklfXHLifobg6ds1Z5v0eTFcvRheDp2T0+LJdOmlBAQAEAKACgEBTOpgFAoKCFIQAEBQAQoKUh0tOzX/O68Xub96PAKD4n5uxz0LPXKsoH2xzh7hx7t/0bMt383w156z5fdsPoceY7eagAgAIAUpAUpAQFM6mAUACggAAIAUEABQAYrk34vl39DfN27uKgHxPz3LpK9mMFlioZDG5GZej8u70rn2dVcpv1YHz+zM9vLn/AEOSkAIAADkCkBQCEAM8mvqAAABSAAFAAIACgwPn9WJ1be/2adl6ealIcTwDHLyvPH6S8CWQ9PwyzJ1+Tq9S58sAuSxvx1Z5Hfr2b1eAAQAhQUoKQpCkIADPJrygCgAAAAoKACEAKSXWPM7cRjnuPpcXe2a6ciHxPzpLpx0MpxmXzuPJd1xu1S9Dh7fUubLU9+Hnm6b/AM2e44Nv9fz+VggIAUFBQQoIAADPJrqgUAAAoBQUFBAQgB8NeeteZ24vK+ger51BQYZfBjCS9eXA5Y8LKer4ZbMukcPd7Hqx7W/T9ezT+etW/wBl83o3L1eDtbMAABAUAoIUEKACmdTXFoBQACkBSgAoIAQAx/NuwfD1Y7bN+9LggKDFr4XL5lljzLjlwyxHo+GXoMvm/F3+54aftu15rt5/LfO9Ls8W7cvW87L9GigAAAAAAAAApnk1xRQAAAAUpQAACFBDX+DrxPLv6/Xr37u4QANeX8/RjVxFx+Uy+eWPKXdpfR5fNeLv9/16eezHOd/LqfB24jj6Nm9DjzvXzUFAAIUgAAKAAUzya4yiClAIAUFKAUgBCgA1nzO3C69uZ7ubZunmoBTWpfGKwuNw5i8nC409Owy9MXxLh9D9B4aPpnjne/lxfPv13z+zO9nLmu3moBQQAEABQUAApnrNcmRIUABYlKUAoAIAAU+OOWs+X245luXp8PazwoKDXpfCF0LLGnPHP55YU9Ewy9YPE+D0vdpo72WGY7uf4a8tV8rvy/Xz7B6HIABQQAhQUFAKCAz1mBlAlSAAKCgULEAABQdHRtwXD09C3efU4KCghrcv59O1jlrGeHGZfPLHlLuMvsceN8Po+yzTlssMj2aPtlNQ8f0Mjv07F6XGIUFBAAAUoKAADOWf/8QANRAAAAUDAgMHAwMFAQEBAAAAAQIDBAUABhIRQBATMhQhIiMxM1AHFSAkQWAlMDQ1QhY2Q//aAAgBAQABBQL48RoD0A67YnR8eNCXWihtidHxo0I16iUtabYnR8aNaUBaANuTo+O0rTcE6Pkx2hOj5TTgGxJ0fK6VpsSdH8HJ0fwcnR/BydH8HJ0fwcnR/BydH8HJ0fwcnRWta/wUnQNGoOAfwMnQNY1pWlab5VYiJXV3RTSnH1HakFT6kqjQ/USQ1D6ivgpH6kqBSP1FYHpncsa/oB13hOjT4CVuJjDg++oD12YsJMzZoezEXjdza8ewSJDM06QaJ9ukW6aTEsAzUbvLYYLSTuwhCm5peJqM+opgqNl2ssluSdG+evkI5CbvdzInhLWPLAtDpwlAuiCKcynGystPmdMC3A4USLLOCPpGTcnZpXA4AI+fMWSfXCiduxZJtmUvCoSsi8gpCBWgr/zMQ5VSbcnRvZ24G8E3eOn9xubdg2bVB6IQjt3cXa0e3nbFXks1FJZc5e2LgXnHERXUGivly0jInSosiRRb7sdFC3ppJJOQei7qUsshkYa4nttOGD9GTa7YnRvLinkoJmQribeQzNqi1k3gQLiSf9oSNJq4iOo6d1DX/IetDoFadxTCWm8poSFkVY5QJgZRKRtVJdtEyzu1ZFi9SkGu1J0bt++SjWj58vPycIwbIs5xUIcHkiRJI6hlRMGIj3lDgNftxGgDgi5OjURJHYuSyqkmnOWzm2s+4xiHYd+1J0bu+50Xj20YdNNpLpliSO5PwepjF0r1L/aDuD1pNUzc8TK/bKO7XfBckMaOVsma+5xm0J0bqdkwiYuBYjLSn2js4PZPN2suLhcS92vd/c1xKBRGmymhrclDNySnNlkLYkBiJ3aE6N19SHvhtqKV7DJyKzFpJK4gAEUr0/PStPzE2oYCARzkuZ3xDITwF+424+GRhdmn0bq9nAr3FHOVmTeYkTLrCoVRQ5QLXr+Gla1rwSDNRylyTdw/iHdWgnFlrlGnarNbtBJRH6dueZFbNPo3UwqC9ws5EpiXCImWAqZw9PwwxL+EYTN7PE5bqtaH8NRpiUSvINuqdrcrAiLD6am2hOjdSQaXECLPlTAoaGIXTXiHdSjbWP8AwgC5SVz9z/8ALXSk8gUiEzmJcJVyMvpqQeZsydG6uxuLa4YdoCrOeRVTE6eIa8TU3T5sEcMT8bYLrJXX/s+IhoHFEdVot2bk3JIGWT+nCOMdsydG6+orQU5G3VFl2cymogY6WHEKGoQObAvyYPONpBrIXX/t+DdPmqu0+X+DXQ6jJ0VBGedA6kbVZdhgtmTo3V5xv3CDgH4sncuZZZq7Jkr3130FD62qOcVOEwkuNnh+susdZnhDoZ1KG/U8Y9mVenTlskzg440zLlKBC7MnRuhDILmiTQcuzm+1tZM5FAEohxUTxCyxySudPF9xswP1F0D/AFrhDocuPeKc1zwao89SKjG4HuBZPn2FDCzZ7QnRu7ngizkfGPTxD2ReoO0XKJlDcDoZx1ljo7u5LE/Gyw8Vzf7qgDIVw7FHcWMai4PJ8qNaWzCHnZIpQIXaE6N5edqi9qFl+xHkVzSYuWh2o1EpA6h7OPjLXglq242WHhuYP61UShz5C41OXH8I1NEyr5BrGIsGTq4H8VFoxDPak6N7ddmdoNHSisYqco3ApIMjMl7RNqWGJ2W6LsJrHa8AqzO5G6P9xrVrJauLrV1UABMLZqLJeWes8YqIdzzmHhm8K12xOjfXFaDeZp5HvoB0yeoqO4XkEmXifZruuQmcZwCrRMJW90F/qVWs3wZS5O2zLpEkWu+l1n1QFkOJAzJkjHobcnRv3TNF6jLfTwhqj417ETU8YGkhJiRRJ03SSPQVZ3+Fc7XnHVbIpHYkBrFOHSjxzGWRIyFQ1osofdE6PgTlyK/j0pFZ2iApyluuYjgFWgH9PfsivUWVtHKqijz3LOLaMA3ZOj4KU/TrOh1qQlzGLQVZ4axmGRjlqITze7wnR8FJNgXO4DybiZJovNeFnB/SsdBx1qFJ4d4To+Cflpx7NwNFe3UFWeH9JoA74omDHeE6PgnYakc9yF0NTFZUHpaZBJE6a16FaFxbbwnR8E59pwXJG7zqg1otJeggc5BNkkl3J7wnR8Ev7Zqu0RLJ6UQO9NQBEO+gAcSdO8J0fBOPaOpV0iAytJeqSIFFEMSHMGCXt7wnR8E59vklq4C4ydIdYdRD5CuU+LcdW+8T6Pgnx8Ev+p0+clTb3g6yeXRRpv7G8J0fBPigcpx8U0OslTT/ACP+6IkUlNv8feE6Pgno9zgdE5UdZGmvcuHWFB6NP8beJ9HwTr1fGxbXIQicvSI6HDrKcMy0y/xd4To+Cc+5JH0aTXJ+5UA6AkOtKdx0T+JgOrXeE6Pglx8y4lOXHcB6GamSIj5hE8VGHs7xPo+CWGrxWwbcP+Ig2cYqXxgOlRw928T6PgR7gU9JSOLMOnJCpr0PTbZ84NXuOOhqj/CpvE+j4FUdEzD5rdwcoOREzhTDMei0DZwTodB9KZjotvE+j4FyPgfKYNXF0OItwYcx0oemz1x+1HVE1M5g6k0zP4t4n0fAuzgBpRx+lk0uS6rWjeligChVy5pKsnLKUTNoO8T6PgXpeYa6jC3DibpsM+j71SkkBcW6xydM2p+Y23aft/AGHEqviM0ZIyb+aboMkx4D6WUfGaKHhRS5sfAm/Ss/Y3afR8A5HRI5gIa3CCDO6RcLKNF0266ggZQfS1j8udJUaT9RD+U4ZDvE+j4B0NPj4so1LksbrWAjcqZlTD6j6QynKlS9x2hwReaAjJsjedu0+j4B0bxSWpgANAuhkHJbPFmSpzCcxvRA2C+vmSsqSJeFMk5K0N527T9v4BcdaIHOm6vB4gVvHxi0mYxRKY3prTZXNGbhPvdLEkLZdMj5o7tP29+qOJPU8KHNdVdDdJvCAcxDCOom9KiXOsYioAurwZA6Sjx/p5RyLuk/b37sfLMfl1BJctjV0OQcsoyMI/IYuBjelW2mZWIBPFecTzYxZvKajqhuk/b37xXFV+tiyZJ8trV3nIWJ/ejcLaEP/Opm1CUDKOZrAC0YpzG+6T9vfuQAyj9oB3HoCigJJ3MsdwxjGDV02ENDG4WWIfby9yKheaiyLgsx7lN0n7e+OOJTjlTUOfNUb0vD/XcDcLEN5iXtoGA6KheW7a9y+6T9vfOjaJB7kAGfB84K1aXGC+McxQct/wBzcLFZCUyXo3VFMXXiVQP5u6T9vfOu+nKnLbQyXLY09NgzvUTc+v3NwtEQKzIHfOyq8RLspttKJoD5e6T9vfOD+ZIj+mQJykanHJWkVdQrjItoQikR+5uFttuS3DuO4iGssS4LcVgjQRxUiEjZJ7lP298ofWlw50pwmjYxd7nE82AiFfubhFnBKEEfG2965mwOY+ILy27QfI3KfRvVjYph1R4c6X4XC6K1jLjXVcS/2JYsWAUetaQbqkgAHMEPfkSZsmXhOxPqXcp+3vXx9E8sRt8nk8JoE+zXWpzZ4Hq4I/ubg2xG2GK+TAiuiyxc0mw+cz8Km5T9veux1WemxYxifLZcJ1crZtMOheyYMFuy8vEh+DLtf2WCE68SqXDhjyl246ONyn7e9XN4358ykLgThMNUlnU6YFJdWfXeNCIHMJkPAdqACwfoN4i1DcyEN0B3hIKYuW58T7lP294buKoJsPEvNelFVKcNRqTxOv2RWYkE7beLUSzzpLfY45sTssS+OjZSwDDxv2lt/wDm1cFVTkW/64G5CJB3huE/b3i46JiHmRqPMkFz40LlJumvcbJGnF1tjmLLvzhypt3QWuqsKNrM06bMEGtGMBASdpOFij4UTBSphOKI6kbjqjuE/b3jw4hRR8TMOzkmWjl+clplMKNtskqTYIpUosg2pa5o1Cl74blpe9nR6XuR+vSrs6w2Op+tJ6XC/cRcxG3M3e0j7jMfJ3Cft7xwPnAcCEWmGTel7wYJ0vfNLXjIKUvNvHFAYyykrDHiUDHKICPAAqzlsZsvrdSJBcrpgmNmuDq0yHcp+3uxpdTuvNU3KOU6YicayHiHdS8k4dBQUFCOtWyfCcDrvTwtwUzPbqPZXTQdF9wn7e7WNimYdRklQ/8AQ3U+NI1qNahWlD+cMUQk/Q96J5xJKY+6gOi+4T9vdvB8AeJeTd6LrOAUA/45iBeLNymgQ0iUznXUbmT5kMzbHduFWgMTAbcp+3u3Y5KKqclrNN1SiOQVkNZDWv8AZaqcxnKJ82PsON5rmWJ56Y5IJmyJt0/b3a5/HJmxYNGxBj5WxkXFSMO5jVBKIf2oU/MhVQyTh48sZHy5PE0HVFoOrfbp+3ujjoVQfDJea7DuClUSLklbGRWqQiHMapp+WPcA4jbKwrQXqRHvSlC6ptO4GI+Dbp+3unRsUtNToB2id/BZBNwnOxSDdvwCh4Abw6a1Zh8oYnS1HVCQDVsh3KMh83bp+3ung0T3Lf8ANW/BYDilPxwIw0c0B66mGqTR2FDwSYrrJuIZw0aWMb9MQe5JQyKp3IKIgGh2w6Odun7e6cm1WXPymUAjy2X4D3BcxlDQeolE6oqUHrX7xRsoSeDKAsgfMTp4+SZPAEBBTupM2im3T9vcjShtakx0asU+U0/BQcSXLIoOI1kRroqmYo6YmrSo1RFvGvF27i3LQHR0mYSjcMYtJJNJN3FKNLkbOyFPmiA6htk/b3KxsUzd4PQ5z70/GYbg6jboZg0aW6Rmo/lV+0KB3DX7xn/z8gTK3rZESu2yYp0kAleyMO1lCzcQaLk2KxVGbY2SG2T9vcvB8AmAFWX6iZ/GUMJI29EhRN6DmOJeH7xCpBiFi5QVvji7HuOTuWq5m2UnHacqMPm32yft7mRNqYFAEbZ1UN+NwOCt4i534vnke5btUFm6iJi8Yt8YsRHuCuoqKNgc/r6GqdQ5lItiKHjS8odsn7e5X8S7pAhGdvoclj+NwN01o2/dPvdtKNyO3qhnBg4fvFoETgGJcmTIdCa5EHp/aRLq3QHRRqPn7ZP29wqbBMxtSyZtEmqfLb/jPAYY68ycuZ9B9aL6V/1FKh9ohRFRJoHc1NmwHoTHVN0GTcncdLuW2yft41jWNY1jWNY1jWNY1jWNY1jWNY1jWNY1jWNY1jWNPAHkglTtAVpDGsaxrGsaxqeHBpPrjKyjfBjEJsDqKlaGrspq7IamTlNGMt8wLUi3Eq0WQRiwTESty+UYmpeWIVgNY1jWNY1jWNY1jWNY1jWNY1jWNY1jWNY1jWNY0mHg/8QAKhEAAgEDAwQCAwACAwAAAAAAAAECAxARITEyEiBBUCJgBDBRE2FAcaD/2gAIAQMBAT8B/wDJvj6Hi+bZM2wY97i+DpMIxqNHSjBjF8e5xdRs5I62dTMsyzrYpnUmNGLY9ul2df8AP1ZFP+mPdNpDebr9Sli+/tdzKVmv3J4MWfslZPBnLMeUZ8ftzgwJ+B+zVpM0Zt+/Pgwbqz9kjTyNY27cGTJkjq8FRdD79ZC/ln7P4s27OnCz20eZX5Wz2/6EmrP2X/Y0vHYhrMO2hyK/K67dbP2WMjjjbsZDWA9+yhyK3Lsa7NbP2KMZHHF0Mo8SpyfZQ3KvK9OPVIqrHZmz9irOJrdlHYq8uyj5KvK/4y3ZXfy7F7RGMmLyjgosr8uyj5KvK9FYplR5ldWfs1Zq7WaeSmV/HZR8lTlZakvjDtftU7NYtT1p4Ke5VWV2UdmVORgpRzNH5DxG6Rn26ZoNFH+C0mT4mb0diryt+NHXJ+Q/Fkhv3SkU1qSXzRLj2UV8SuvlaksQKuszYz7yD1JPBjQxZFLiVo5wxR1EsYJSy/fIlrHItbopcCUepYKdFp6lR4g39Ah8okSW9kU+BkRXfxx9ApSwiO5PlePC9d6pfQKRHcqcrIjxV6rzP6BDcjuVeV1xV5cn9AhuR3KjzKyPBpZ7/QI72qWRjS38Hv8AQIbiRV3sjqGIe/0CG5kq8rI8DQmS3f0Cksu1XlZHg3tLf6BS0tV5Oy7Jcn9ApiJ8nZHi8+T+gUyO6Jb2R4MWqcn9AhsR3HbweBbDRV5fQIbC8u/gXE8DehV5fQIktIO/gjsR2tW3X0BFTglfwQ2I2rbL38dzwVt8X8FPYharx9/DcS1SK3O72KWokRlmWCotH7+mhLDyN3exSYtxZjMa09/T0WCUvg32PYp7nk3mjONCSxJ++RV0gl2MhvZ6TiyqsMqcvew3PBWeuOxkd7VfDKusUyr72BHkio8yfYyO54KkeqKwb0kVVp72C0I6Zd84s7eDq0FLQqL4v3sSWlPtdlsS0iRn/CWufeLV2q6RS7XaCzEmvifixUpalRYkP3cNz+IrP5XxZ2py+OCT+LTPxnioVt8k18vdwWhFfIm8t9rtTJIovFRFRaFZYl7uO2CMtG+zFnamPcWjKmsclXx7pCJaU+52gPcloxPqgVOPuobngreF2JWdojJx6inpHBNaP3UBbpFV5l3O0dxmSDJ7+6itCPIer7MWlZb2n4IyyPPkej9ykLSLfe7Lc8FTY/H5lXcny9xHV2npBK6tgRKytPYpPE0VCqtfcU1ratvjtyIdluRWhKOjIvDRPYq7e4p7C5FR5l24Eh2WjIy0M+Lcok18fcR2SI6ZY+1MSY0YMEb0VmCZUWj9wh6Qb7EhRbOk6ddDpOhCwjB5JxaZRl8MDevt47ngqPEEhLJ0M/xijg6TRGUdQ5O3gYyOhIlv7amrT+RDEUdSOs6n2ZMnUhPIxiY9ipy9tDYfbk6hs6huyQnraCUtycekTyir49tFDMs6mZ7M2VmyO9urpR15ZKOIlTb2sVl2jDqRKl0R0M2x+iEW7S4kf6PWJNfH2tPc8CkoJEppkh/oRGeFZ7GxTeYjXtaex5wVNXgeUZZkz+lbWkyg/iPce/tIrQjyJvMmxS/poxr9UdhD3Px3oT3KnL2a3ER2b7Oown34NiLzaW5Q3JlXf2cFl2lpT/Srp6WgMnuUX8yWxV29nT/o9iu9Eu9LJJC7YjJLqRGGHm018fZwWh5K7zL9Ge7xkZnSyJbP2aRDkTeZP9K7ER4jQ8Le0Xr7OOrtHSLf6ESF2LcjxJPJN/EUmiOZ7DTRPSXsae54J/Gn+pDv5I8LS2t+LsTKyxL2NJH+j8jZL9CsuzyQ49n4z3RJlbXD9jHSOBPLwV3mXcrRJC7PJDbsov5EifH2CWXaG5N5ee/xdW828lPYe9nuU+SGS29hT5GRPEW/07LvgyXI8kt7Z/5P/8QAKhEAAQMCBQQDAQEBAQEAAAAAAQACEQMQICExMlAEEiJBMFFgE0JAYaD/2gAIAQIBAT8B/wDl6lTeLyVKnnZvK7lJU5IFdxUqbSp5mbly1QYV/MLsaoCgLsCLF2kIKbTHLkxfOV2D38UIs+lNtFryhyuASUBHyloN5jlCbAEn/gIm45I2IQEBSv8A35dVKcPaHJmzR7WY/wCGVoYsOSKz9IGdfhdkEw9wx6I/dhyeYwzOGqYYun2/ATYcmCfeEO8yMPUbF0234MrDkSpQM4An5VChpg6naun2/BlYcibAzhrb1T2jB1O1UNl3mAqZnBFhyLrA4Auo3KiZZg6nQKhsv1DtAqA8cB5QhAwpuDK6kaLp9uDqfSobL13TUTBDbmw5M2BuDFSFX0C6b2MHU+lR2WOSb51MBQ5Uj3YGbVcqkqttXTnyODqdQqOy1Z3awrphL5ueYIlZhArqfRTj3UlR34Op3BUNlurd4gLpRkTYmUBzRaq21MM0iFTyeMHU7l05lluoMvVDxprVARzlQS1UxIIQycCgb9RuXTuiQpKce4lNbA54qnk+ERBwdRvTHdjpVSuO3JUh3PH4B/jUTz7TdBesPO/TDyn8BWb5JypHwF6ub7ELphAJ/AV/tO0VHYL1N5vREMH4CtonaKjsu/ebsHiPwFTanZhURDYsUd1pTdPwFTbalmLFTncafgKm1EqhtsVGaARTdPwFXaoGio7bFe7ESm6fgK5htqOyzl7uzaPwFfRe1R2CxXu7No/AV7U9gsV7vT2D8BWX2mbRYr/V6WwfgKu5ek2/+kdUCqBmmPwFTch6GB2T0dUFQ2fgHnMqnvF/aqbk7W3THI8+U5Ut5wVdydqsiumyJHPv0XtUNCb+1X1T7dOfLn6ui+yqGy4XUJyfT7WByomHDn6xzhDMIADK4VcI6Iw6nCaYPP1cySqbfIDDW0XpM2IjNMMtHOnJOVHN5KOCrttTzYU0yqOznauTV7VAZThqbUFQ9hDIldOciOdqn0vRKpiGjC7Re1SeGOIKdlUMLpznztQ5qJgXibnRaFBndmnNgqgfMc69MzqAXmws7cqe6E6mHapvieccYFqIlxOEWqGHqkfNdQ4tbkmmQhpzdXRD2VQHjNybC1ZvlKYIeIXVCaapHKFTMsHN1XZwifFMENGEWr6ph0KqiWFM1XTnw5t+pKjMDATYWroaI5tTdyoexzRyCJlMzqYhasm6JhloThFQqju5qoYavaoDMnATYWq6JqY8s0VUy7uVI+Q5qr9L7KoiGYhapogmMDgqlMtVP0eaqHyR2pogXCmws7Re1R9ohGATCaZE8yTMqJcBgFxY6I6qjuK6jJiYZVLNnMPMBDVU86k4ZsLFHVUtyrCaZTF05kcxWOSGq6canDFhYp5zTHeQThLSm6rp8iRzFU5wv8qkIZhlShYqo3NRnNj4vVE+fMPOZKJyAQyGAIhEhAqVKqar0vSriKhVI+Q5c6Iym5vAwEwi8NX9F/SQu8ovcEXyi/uK/wAqnUDgupHmm/fLv2qM1REvJTjC/oF/Q+kZJzUj2V3BSfpeRUW9oaIGE8l2qYmGW8tWKn2qZ7AnuJKlyg/a7Au1dhXYv5rsXaqgQTGhwT6ZCGqonw5apuQt2ldi7F2qEM1Fyqg8UECRomO7tVVABkKgdRyzjqqQtAUYIwQqm1DVMEuXbARf3FUN3KvMCxf2aKnVLzn8dRwhe1S3py0cqR8xytY5QvaDe8lNZCHwkJzJR1TMnC1QQ8ppzHK1sym/ao6SslChR8LtV7QXUiHoaJuY5R5klf5VMQwKFKn4qmqKbouqGYKboqRlg5N2QRX0MEKY+GqINm6Lqh4piobeTqmGrVMzqfIbVtUFT2rqM2Juqoank6x9IarpxLicbjATTOCVKqoJri0p1UOaQUFRPnydU+SGkrpx4z8EYqmqC7Sc0URCpmHDkinFHaqYhoGII46uqGSpEyi0HVPpkaIIcjUMNscyBjCcm4quqaFTEPREow3VSFTMtHI1tF7VMTU+I4PSqbl7TN1upMIKgZZyNc5wtV04zJxhGxw1NbDUW6oZApgVD2ORfm6VECVQHjjCcm4qmuDqB4JipHy5BxgLVO0TBDQMYuber1Lt0VUSwoKnuHIVtqhES4D4dThi1QKMl6TNqOaiF9f9H//EAEcQAAEDAQQHAwoCCAQGAwAAAAEAAgMRBBIhcRAiMUBBUWETIDIjQlBSYnKBkbHBBWAUMDNTY6HR8ENzgpIkNER0suGDs/H/2gAIAQEABj8C/I7cvyQ3L8kNy/JDcvyQ3L8kNy/JDcvyQ3L8kNy/JDcvyQ3L8kNy/JDcvyQ3L8kNy/JDcvyQ3L8kNy9B3pHtY3m40Wta2vPKPWXkbNLJ1cbq8nYmj3nr9hBTIrGzQn5rytiafcevKQzR/Iodla46+q43SsMd8bl6B8vMO0/dtxcrljiEIOw+Jy7S0OfnO77Jsssz+RY3ChHBRSCG9SVodfNcDghdskTf/jCtTQxooGfRTyGKPVYSomyWWOoaBW6FFZ44uy1DJIWnhwVbPaK9JAjLZ3y9k1xF5msw0QbboK/xIv6K/ZpRIOI4jem5b+ZbRII2DiV2H4eHQxHC8PG5fpE81GVxAxcrParHHTszSQes0rtS8BlKgq1sYx0sE3lhTCh4q0RsYxoLeGJCYTaaYeayn1U1yWbEN4hPa6Wa67ChcOaqJw73o6q1zTNZK99GYGlAEY4w6OWTVF7+qiijoWsFKjimwQxNaW4yzN25Lt7O9zmt/wASLaM02H8RAbw7dv3QcwhzTsI3huW/XpDelPgiG0p877z2t4N8LAhLF5WQ7ZDtX6Sygil8bOZRZEy41wxrtUjXOayQHxPxTH4yPGBJ2FXRRo+ap2rgOhVb7q5rGRx+K/aEjqjVodXFRnGO6nGGV0deLDh8ke3HZvd56ENj1jJh2irZjSYc9jkYJQXwg60LuGSZPA+/G7+W7ty30vOtM7CNnNGecyPaXeUkHmq7ZgOyG3n8UewPj2Dg3o77IvtD8DxP2CusN32uKqcSidOxY46MFXgsDRXZB8QhKNaopc4U6ckG2dtwuNKecf6Zoj/qNva9U5jgblfKRc+qjnhdejeKjdm5b5JaJTRjBVdpKcXGgHBoQihLXt87rmj2Ty29scw6zP6hEOPbyO+PzVXOLj1VFl+pqdmigxb6pQkYal2x32QayjHu/wANni+J4BGVhvWkYnqv0ed3/CyH/Yee7Ny3z9CjPkYTre05GaQNkkl4baN5LtGAv5NDqPGR+y7Rzr8rvCD5vUrFdP1dFXRgr8XlGP4H7ryTm5RY0zcmy+Jsm3o5djIazwap6jgd1blvc1oPiAo3Pgh2msweUkrxXaxUdTzSaH4OUz5JH3YsAyQ4/NOlftJrRVHyVP1vXR2bneSccU6yCIvDcW4gYJ8DWMIPFuIHxUJcbrS7s5Burct7stlHWQ/ZCeN918h2VpgnCSSRjqbJWAg/6go4MCRrvI4uK9V24U4LHBWeWUmUVuOZ9EC2GQtp+7oE+WMUbJrfHirLM7xFtHZjDdG5b3aBwZRg+SijdE1jWNpVwNPmKqNruxezFxuPrgNqc548RrgtU1H6kBAfqHRB4beFa9RimmaZsslP8V+z4KF8b2G66lGngf8A8UsP7qT67o3Le7S53h7c1+avMjlkHstTpBBdAbRxIpxXFp7te7GEwez36BQmg8Qwcrl9jA3DCOp28ynvvOc4O4q3N90/XdG5b3aP+5P/AJKr2xsNNvhU/ZvkLajjUKrXV7sUnPusyKZ/l/qGuoTQ1RLbO9oLq1E1Eb51K0oXXuOStzvNo0fXdG5b3axzdfHxUUrZLtWjzW/0RDpqtdtqFgb3dhKcOR7mTUP8sfqGdpUMrigY3PoW7HQk/RMiIpV17j91aZPWkp8hujct7gtFNWRl2vUK412qw0u37v2VDBHR4ILqkrbXu05OKmHtdx/uI+4NNEB3KSSdm0BXbrS3ZWJ1f5Jxb4Wi6FZWUo5zb5+O6Ny3uWgrJD5Rv3RbS92gpTqi97JT0ADQPunyNaIwfMHdtDeT/spOtD3JvdUnut+ml7/giOQ7kVfK1FSxpxCe+4w3B4XDFRQ8HOvPPTig0YAbo3Le6HEJwZhE7ykRTaDXIo7oU+MhxfXxOwocu5VWtmRTDzZ3LQegU2TfppaaeLWUjubtNLzWUFalX5K9oPMcuxjrq+LGqdbJBSSfw9G7q3LfCwYTs1oz9kWSgtbW7I08EQMW8XAVKL2sIpt/rpEnIBWhvNlVZ3ZjuWj4K0fD6aABtKPsM7gBeQ3YHesg1sjzJ5oJQLwTAw3pXc+iAAoBw3VuW+ut1kb5YDyjB53VdjL+yrt5IiCJxbzHFa7aV0SM4i8EWniwqN3J/ctGYVo+H00Qt5G8rvFxA03Zth48kS17w92xoO1MibV7uLjsaEyzwjAbTzO7Ny359ssLfKbXwjj1CuO8HFh4IuaWsibw4rsziFaI+ocgz2nNUh9VwPcn95TZDRJLTYKKKPNyoBUpj7VEez58lchja+T1+SbHECQPFI7Y0IQwDHznna47u3LfzLGewtXrcHZqkrXQu4PGwoyWupPDkpBZ/wBk5nwqrO7g9zSrT7te5JhXWV71m6C+m0kosL7gwbUqN8MoceXFXBqM9UcU2W1g2ez7aec5NhgjEcY4DeG5egDFPG2Vh4ORf+Hy3D+6k2fNWf8ASYHxi9dvcPmrFOYw+puY8MU9h8L2EJ3ZziQClOul59tRvrShIJUg7XtKAXS1Nb7ITy0eN1brQr0jf0WPnJt+SD7vbz/vJPtvTcvQRChhnvXe02tyVylcKYomUxkUrqu4aSfbKljOFUx0sjbvFo2qGB+Mch2BUs9nji6gY743L0Hf9U1+Rqq9Vb7NaAZJXODWycg07NP+op3ArHaAqn/DZvrcvQZa/Fh0PlZO1xcdaOuIOluZR0TSc3U31uXoNpRU1ouHsLwbf4VppZmfroKZ1x31uXoMZopk5eS101A2uA1dMYIIz0PPRRD2RvrcvQZVBzUDHOHZiR1Ggceuke6EbjvOUmSblvrcvQZTc09ocbpJdTrs0DNZBYKWoQy31uXoMplMcU88x9zoGaNdYniVQ7U8Vxom5b63L0IwEVUmhvvBHRI4EUuqM+yN9bl6EbkpcKbNEfvhFEP2VwcpB0UfujfW5eg21xWTVN8Ppoi98J2h93io/dG+ty9BhTHkxWj3tEXvhORRUXu763L0GFaD0opmspTV2c6aGe9ocONdEeW+ty9CO9p4U/6O8SRVwcOOGgZoe6FJe2VwVE3fW5egz0Qyc7+X/vuQHnE1OV4H4I9HHfW5eg5EW+wB8z/60hWJ3OIIkLFSD2t9bl6DHUp7JJTHGJWtJGSkaypYHECu3QFYj0p/NDRIOgO+ty9BFDk0VUBii7W0TTF7QdnhO0/FSF20uNaLydbvtIKL2ZCEzlsXRN6t31uXoKitLhyuj6LsGNY9kXhrwJCqeOgKdo82VMq0tzVrsbqXR4BltUVcDXfW5egh0FVEw6l59STyCdS0std7HtGaQrY040uuCCP4m4AWf9KLNuK90763L0FITspdFFdvE0j+vcCtLOcf30WwbTHab381FJfpejxFOKidzaN8bl6BJTBzNVanTxtljaaAOxCtXY2Vgu2V3haBTSEB60bgivxWLqT/ACVz1SgOWG+Ny9AlOcdjGp0h2vdVW8NrHDFZxX29qD5YG2hnqOKcWi60nAckFZOpI/kiraz1qH+SlYnjrvjcvQLQpj6+qoW+zVfievQ9lG27zxKusaXu5NGmxu/it+qcpXO44J1NhcU7q3fG5egXHkFZYR57/wC/qqL8UtErg94LGsrw2bFfheWOV47ToidycDoj7UHspRtHBCaJzXjg5qjPMU3xuXoE9SmDhG3+/tot0N//AIh8zcByuhSCG7qNvG8aIgihGmzv9ZgUcfadm9tS0q46sZPxa9WeTndO+Ny9AFM+atU3Wn9/LRarjAK2zbx2KrSQeix26bCf4YxUSsr6eBxCYOQogd7bl6ApzVol4NGCB4uOh1xr3x/pTvLeZxwHNTudaGQmNtQ07XItO0YabI9xFxtRT4qBzW+cj0cCnM5FMy3tuXoBg+KOt+0fRRN9nRZ420/5iQ0HDE92Km0V+pTHdVP7tUa6reaPR1N7bl6Akf0uqyQRjjU46HPdg1oqSrE/sezgvP7Nx8T8dqtD5rSI5GjUj59VTTaGXq8ctv8ARc6BObwcE0dFKOdDvbct/JTRzKceEY/v66Cvwgfwyfp3bXHzaDoYduCPR5Wbd7blv5Q6BTzes7RLK7wtbwFVYHTsuVhFwVqaK0Plmax4AutOfcntJNKi6G8/7oinXTsKc/ZU1UXy3tuW/tarQ8baYJnXRO7kw/RWIObdpAKDuBDVodXHn405Vjxje0EsOwq6Dcl/duTTyO9ty393QKNnrvTG8hotL3eoWjDimutDDG8xjVJqQE+2Onbe2NYDsz7kdo7WSt+PVvauLnBFPjtEd6mxw2hMe1/aQuNGu4qIu8VMU08xvTct/f1Ks8XBor/fy02jjq0RvC7RjcO6XioIfCT/ALzodkhUeF4KLORTemG9Ny35xTR8VPJ6uA0vJIBJaAOeKnfMHNcaUDtoFF+mP1Wu8A5oHTNMLQbnk/J0w8RUTuYQyUo6VTgnjkd6blvwHNPdwaE+Q7XHTG54GrKyhPDWCtTqEYjbkuy7R3Z1rd7lpo6p8nhX23Kxmn+G36KNPbzCGSeOeO9Ny35g5YqU8X6qj646YXvoGiZhqc1aZnU1n8EbRd8nzPFMfwdXTKBGx8Duz86hGuVY3EUY0UzQeBsPDRTk5N6jem5b9K/bQUVniHE3kG8hp/D3SC9SXicNhOz4K2Obi0yuUVmkja5seGqNoWymZV8uqPZxWF4at6rkYpX1JMerTk8kpo9V7h/PTM0jY5Qmtdam9Ny30q80XrzuChZSgbTb89FWm8Oi2fNWMPIIa8uI/wBJVoMNwVc51adVA1zX3am87ZROPasZFQgOdidipP8AiHwjIC7CzF/bOF2/iUQ6aMMT4L/aVN6tNDeB5FOfzaFeYNYYjHem5b8ByU0/LYmoCoY0ZALGdnw1lqRSTnZg1Us34eI29VrTCEH1VW0WuR/xWLb+a8nG1uQVXEAdU5sbxIRtumtNDgDsKBJrREJmW8ty30AJx4rqUzsrSYWjAhqrNPJLmV+yBzWqwBeUkZH7xov+YDzyYKryUD5PeNF5OKOP+axtTmjkzBa8jn+8aqdvOP76BJC+gcwVadhQZL5CXrsKcqcjvLct9ceQWsQ2vNa9qjH+papfKfZavI2X/e5apjiHstXlLVIRyvINFXucaBNMp8qaYDYmXdtNbPuNb6zCEVC54rqkLA1Cma9znXaXalSD47y3LfX5qyWdlS55rQKjmlp5HvMEspkuC6K8u7ZOrqfyRUL+TqIV5qnrNRHNu8ty3wlMCikOyCm35qM0bqch+rszvVkGivquBVVA/mozzw3luW+U5rIJz/3jyVt713h3JL8Ikcbt11fDihK0FtHk0/1Jp5q0DpVRQM8TzdCbG3ZHQJp5HeW5b4ByU8vJpUTrjhHdwfTD9bZn82D6K0N5sKktjxqx6rc07qKoZJp5jeG5b48oM9dwCjiewOaW4ghF9jd2D/UPhV20RFnJ3A/q7G72AiFFA3hiTzKaeiCb0w3huW9krqSrLCM/sqaCyRoe08HBF9id2L/Ud4VdtERj68D+piccTU/XQ3JNPVEJw5O3huW9lNCPJmHdLJGB7DwcE60wBzR27mU83adneI0Pb6sh0NR6Ip46V3huW9gIk8FPNz+/df2ZAkpql2yqgtMkjpLQ+dwOOqMTsCbGXhgP80+OLENNMO46RsTiwUq740RtEjQ1gkMRxxqrUz2gdD6GmKe12BogU3qKbw3Le8lM/jRV9Y96wXqNYXuIHFVGBRvYmta9y0tvNNI48OP7Qq19Lc5Tt5tBRTWzPDBJ4SVUY6Iz13huW9uUbPWcom+z3XHkF+GWeKQPfGyr6cMFI+0l2qNWNvnFYtuB2IVDptV5r70jGeYaePmvxFsLvDab93pVZsK5jJM7FnaOYSacVdBNBtjersnkJOuxBwNd4blvRQHNQRcvv3rQxxcBcJ1TRfhey8YtjW0HBUtlaebyr1RDfDeoK7e5aP8AKj/+xy/F/wDuHfUKG7SpqMU68bxTKDVINVSaPW4PG0I2dpvtpea5R1ON0VTD03duW9UQanu81v271qI29k76Kwtc8vd2PHRSuFa9y2sBdeETK44ftF+ND+K/7KzH+JoZogk4FlFRY+a4jd25b0xvVPeeCmkPetRc4CrCBUqIm/qsprtu/IKUugE9rcaR3sQEO0F2v9/fuW+LsXvbdaL7B4dbivxmPyl6r3eUZTgmHlIEEw9dED/VKxqCOINFKwbK1G7ty3ov5KV9NYim1bKFx7z77A4tpdrwNU2n7ofdSduy8675M8im1O0/Ydy3PaNZ0LCf95X4uOcr/wDxCd0KY7TkdGY3duW8uKPOqiZzNVG3kO8WtwLnsGPvBOBeZHXRUu71uaIqUgbr89dfid5paTM7D/SFIoD7A0NyT8kFGd3blvTVEzgB9+/GeHbMr81LaGi411AAVhBG+0yuI7R4rdCay8BU0W0LaFtCtEPZ+UfEGXh7xKtxGwzVxyCmGG1Q5aGohBA8ju7cl//EACsQAAIBAgQFBAMBAQEAAAAAAAERACExQVFhoRAgMEBxgZGxwdHh8FDxYP/aAAgBAQABPyHlfYroDquPgTFRJrEmIDHH2e0d2eyMcJhCAKGAg7XbP8xQjiEYZ3AuuObbIP8ABPTMHgVxDyvsNs6b6bjj6B6ghhHEHA8XH2O2dqeR8R1j0zhPAdhtnSPTPOOoIukYaxoeAdhtnYDoqLgOgeyPAXYbZ2A/xRyLr7ZyOPuHzrgOxfY7Z/4jbOLj7Mcx6z7xzbOZ9iOB7B877jbOUcr5xByjkXKeR9Y9k+TbODj4vmfUf+QeB5ts4uOOPpj/AF9sjh4D4CLsH267rbIUI4QeIDoL/KcfX2yVQByACLvCcRXECMAC4B+ELQFyH5R9ozD9Qo0LJ+2DPgv3F3mSD5EWA/iQA/MvAf0gwYgkAOI4PutsglLgIB3hyxgrnph6w1PxIb9QPSHGD2/SEzyyMDJFqxCuakYnoxEcvXlRQIQlS78QnkqJGkIDklUaZ3h6gAo9F1L/ABARXYfZH4l7cFLCtMvSFcnmgfUp6F8fMO62yKERQduOTFG830GcPzMof+Mq8RghpdXlFr5sG4ZztAk2tCv4xZRi0Fq7NR2ADMqVdhlCA6BpP7DCElbDdTosYU6QRF0aQOQAl8gKLoOeOA6Y5weH2AgH7IeNNWcx94aMxGoB8i/MvLAHDwIInBoAh6PsQY1WWwRwPAcV2O2cii6z6dOL1H/EQCtfIPRiE1FoaNFhGfrFj9pw18wB0SCNhG0BHTKqOoEGCQmgsGAwlkFSX2gECFsEQtBMzQCgWROAlplQhlDJsP1CzTXo/wC0gDQhjv494A8c3AZDT9mCzBYG4HgXOHmApYtXq/USFoT7zw+IOMBhcsjkYugouCi6W2d0eKW/OLM6CCtISaHAQJMUM4/zGCtCNuMvBmvhAUpUiv1SxGKIKxDGISXJgZgUwgTDtiojKtg4SExM1iigitwEgZ0rTGMTSijhdmgLECvNEqDWDjtHi2MOgOHjsaYBm9IRhAM+TIdIUGpHNBya6wCZwZaHXrLnc2yOPuqx/muQELjfhpiD00Yalin0Yo6Bekp+I2gHlXU1DMpSqCZQpSuMoSqAWUEv88LpggxmMNSZYBBWHwASRl7EJyXCH6xlF9g2es2PeMfxgwochHKBYv8AkM4QAEFg4jtdsjj7omWth/lQZA0T/wCpj7QNYCjR+GeNUKL5sd9jSAhhlE1MJ5rGE0DcQGWhvDMJgeLhNBki53ASpZkw1Jo2OMYQ021eRROdWWHXoPADgHlsv/F/zEFCWX/kHa7ZyvtkbUbmcFIHSTUsfJhZSVP+kVHgsQZ0gr7WAEFAC0Cg8QZw+OSCcUhEOcwmEwmEw5DBSC7GeJxMA9ACm2hjpmHRfMnIzO/9JuBtHs8YSE2mRpsY+yPDbOV9sotcg7faAl5Y1nAkCo9bg3hFOo8RU7wzWps7nYIe8Gr0sDASZHvCPaX8zSDgAY0bieFpeEAPohceIZwIWJH1FsIu/qAgxKEL1KjMM8GxrX1hAnvYfHabJ3ZMFhEyoPyTAZvK9CBsNYGTCukDwDCJEtI0pw6CwxhOO+ctFiJeaogtGjM1TMZguHwCFyE7xgbXm3kKiWt4krFkgj7AvEc8RAaFP7nH8alI8A/kHpPi4+VQPadEdB9Fwg6IRaBIb3AeaKwqVeYi9BlCHIm0qZG0Tt7R4GDSEqGEvkoS6mBBhfueAzQFxUCIO1sTKF0lAJFhXX8KAmME+oFhSeK4RdltnSfYiGIoKECEWhNQL3CiEUPDq9Z7OqjWNYgbSovAQmJD+Li+CdkSClo+TxBwh4jAvLTghSM8kUUR8ylaV6nVk0M/dpdo2zsF09ZWeDhnZVzzQVrqcwg+BCRpbxAiPppqrKeIPLhQWQlbkTX0HIV6bfqUDy+Q8bzDJXxFGBAMkdOTrAF1AgsaxbTiQAp4AYwx8JYH+M+V9fbOyXRGO8tR+CJXuKMLBrgRxheiYmgkK5rCWuxUZyj0iOXRzcpu/uYGouRqy+whsOXFMAMKzIxInrKSmUE4BwyGzlBEgQADpkcXzCqMT5DuTGf7g6vxwcfRfQ2zmfWXMow+uKn4ODgtXY+4AmigILB1JVUEcFYIwDjKM+BnwhHcY7J4I2ORxNPzPAAcT6rIIwewhPSUygOkKEpEpsaA+4albkENgCDrDjFosBr/ADWCBSQGQ7TbOo+muQZQAgRBxjwzUcA7ehiG+sAT6AqYNjGGPEQMsIkGLWUGsIHAZ/F1DNC7YnkahYHzHaHwOLyqdpkOQiVj0jBARlPQax+CFh+4zgAnIVESQ4AOLbgATf8Ab2im2dg+opFvV/Qw/hIFSGPpEGWGh4GHkxBEYThcpTNx5CL4VIPxMvx+w/uKT+1yVvx+Yb0vr4HqoiEyXTHoPzGzW8WUDJA+ZZQMmhetvHzBG6UdVd9FpHUiX+GYIMEgGA7XbO9GNKRWjBrKwoqCx6wtNhENPOAQNhAyptLhPyI+YTAHXsYusce4/UNIYJX/AO0YjXfZAIpg6j0rCnb95+o84nALJWNIEHRBT7IXEkAeqZiCQ6t8YntBw2zs3H0jiIFqH5NIWAJdCxRioCLbNZx+KDBEAdqQh7iGM0AG9jP5R6fcrvDwVrT8QK2fwwkoerAMfX/kXeFDb6MGzDWAvBgRYw/KAU1WUHqFz+4shw/lvEzXL12Pb7Z2z6JUJlR7D7igTpfQ4xkKxBvrtDuwxS4EaQon7DQxNxX2kGGhUN+BTm708CGq0SdyIMo9c26UEQYNIqNP5ME0afixGRmPDS6YxN1fjw8yzS0O5z7jbO8fJcxkJzPcGP0flGL1xBm6aJfwkO5C94V+4PSB8TESxfiG/ACxxP4EKtiXMBcfBgevIRROLltSATrjK3tB5nCGAMeuP8Xe8VCWE14Yci7bbOUwdkekAwGxCxAosRBJLdRjADFFOOBqEkU1DBic59EunJLyLoZW3zfs9MYUZJQMwArtA9Ewe6/ebZ1j2pZEfwHrACtiUN9DZqRXsicoiX+KwjUlmEEElclEKDi6n+Pe7Z/hiMoDeIoCAMFisb7B+0ZQWMbSxt4pqxrK2YlrYbwP+97tn+GYgF4L0iILV6gYMqGHQxf9lUArmHAg9gBNYufqe92z/Deso9xEKkkbgFVr9S0uQxtqUCxM1MYicwOaGfF2Y6W2c76K7MHAhrpCIuZwIAyXraeZ94K0/gg4IDQaojxAFY4ICeQ9iuptn+J6xFgwkzSqr2A4PaEVLIHmkxSj2MMXzlfjd7tn+GSgEKjV1gGhFhgznNtjRFAnwQ9AqNvMALTBhM+j45HxfbbZ1B298ZmE6SokOEBuLjwzwEn+ys2wgkYgmJGAVCGZrUbbovqOPn2T/DQHXGHfQhROkEfHAWHP5eF1PMg+8oRMYF3pP4GXKBFyDnfU2zoro27EdCgLiCOYZ4EuyEiE/wCesEhiwwTBKCAFnQT+plxXOuz2zlXXfXMMeYMN+J4yY9qTeGxl8gjSv8pX4Ztnx2Lj6eyd+eQ6ek/tF0ltCIqqhJ9XwMXkHzLvgSodBUMrJ8Qn3v2znfE9kec2AyAlzJJny/qYcA+xQZ955jjFdzJAUAOxQ1StJ4ixue92z/DreSXcvgEIESlk6mYhObCO8toAJACWSHSyHe7J/hvbMqaDet/DGHAv1oPEA9hA2gmOjVPdzbvdk/wiYZWHGY+jAslHQbwlZERRAGj4rFog/aQi5giABTyX5HK+42TovsnHzekYKqakpa/bARcyAdsSE4wG8IDPDxcAtP8ANP7juQyPomduL6uDpnstk7UdWkzGY4j6oxdzBaKE+bwhblRjeJnIMopH3AhlEglhHPxH3EmCwI89O/ZbJ2L530ggTcSANBYXADfi0EmxVJL8uNcSBGxgOjrLoSILhdoYuMl0yUCbAgMFn2Dj5ny7J/hPRUDCOsFxHWScz04HhsZko9eA/M+CCOynh/yYAhQBUUBTUAbdF8HHwfW2DtL9V4YCF5EQcFgOoKPYxS8URXBT2gRqbSV//wCx9R5MZThk/OSqz49DX7h+cO7snzuPhsnK+8MlcoTFWR+ZdJ389XCMUzokCfYN6QfAXKAPtGdQOSyhxav2pS4dYJ4U3RD6noEe4KlLLf3HWPW2T/BZ5XMNySepUpIihetYAFOBq/kg+RM4YwIGhGEtQRSiqQF1KAgEU6f9jGbAjJGsoGUfb/vM+L6L5Xy7J2b6yZIRWywjaBDCgAUomhGw2B4N7wSzgGPmFacRBQqJ/cYYKBGIcedKdZwsPWXNjIis8bP1H2D6ewdwOgTFs86fsI+t+AYSzMQ3ch+IHmqKko1MkQcOAEURlQe/QQRjSEAw1YzLaqoPuaavd/73mwdy+dr0hpr0jIUmHv8ApwzxWVa6vvNZBFHxJlcy1MoA40o3WpNgD6GFgx90H6hs0t6TWAPnPI4+vsX+AtVyhRMalPAmvwPxCUGbRYQKGRfwOEYwN4eEOuNZFiKkdp5NLpqlqIACBRBGM39C+4DNmp5l3NJ7d3sX+AMrYAkYoUAHoufiaGBCGEaiIuEJdApiVsjrKRFQRRVRnzLwgMOCAyD9lYagJEsEChjfb77vYOs4+xKCrQDL31fACQPzAEAQ2rTKARMpilXGKYCo1ldPpoS1ZRkzRuJXHaEMqwY1IoFSgCYqSPcQGHhfaKKxbK+uouvsHf6KCHHWTKDWA9vzwUOqFCFVdfGsYx1lEVpX2T+CfzAIQ6iDIbFoEQGwXrDTzx7TYIOK7syyqVWWxoJPn0j5L/HBqbRLC9hDREbolNTgPAgKIhiqUZiSQZlCUwCtYSa74dHIymhQIgEqEF6oomDq8jkfMOx2Dv6uozM7wPI0EyNUfr64BMWL3QocEd7KZvMYDFMUGIMKUzQrzSjTPRhHoZqhVz0zictHfu9i7+oyRjxPwK/iab44HhTQEWQQEI4HF+CeA8CEVSxOefsNIKaoMdoGqjTiBf14aMA6InTeMyl3t0E5GG2JMwxdQxNDw91sEXekoStacxaCIeT+IHBtTFQ80+4f2wg7IGsCEAlG4jbYmUGZQNBFCLzSOohoGYmVXPvR9xK2k4Wrd0319k7l8viSC7rFHzUP6VPzxLvGVSa0Ax8SlUAwLAwLTXOXERJJytApwZNpfMEBJ1CYYMeEt4tapO0NFzISlD+is8+AMEMi+52LmcfVcfR1FqADGLhCO/kfvjfG8N4hekpzSBCjQBBF4UGWAbQFucTCZvDcQgVFeotCGclczog8gSveaqI2l5xSaVAd02LovrPg+XLmpCjsh6lRUybuJ6iMKgE1/SCoAmNBSsL1hFJE5HkNI5IsqDxLpSkGgH/AOGJcqyAEmqEhKAC1xQXqOBRwEE8ph991sXZvi+R8gjpFg3VvelPuDBWAONlOwLVx2GC0AgBFiHLngCDQptFUUGUpIMxQg0RRQf4QSFhSQsCt4CCUqZpVnj5gQ1vkH3L50hpOYgVwQEeobgy5UPdTutij7wnMhH5GCuQjEDHYB5L4hIBkoQFaMaxHW96JyytbIY8wjAAYTU1QYGGIFhisr/2E1SHiCpYsE/AXEBNHoFjSYFsoEu9VhBjTArEqhLrpB8CkIwq1EGAaikeKwCZAygOfc7F032TjWkZbrAGHcPh9RwWBVlhwqcIMKEySSMCJQmolKAg3h0cPxPSfAl7RyDC4nIZ3LpuaIWZlEphT5nqR0uYReJQ1CgPRY36O52KPmcfalaw3UOfDQ50ikkmHwWZpGTUao76oIQ/QSvBhkw5oGKg2teAP3CRV6s428QPjH43mWGrqsPQPzwigiyqUSLSggtEftGYCxDEpbmDudi4uOOPqHp1AWLGUHqoxKAq2MABO0Zgc0BupeHqfWINI8wDu46bsBAewgFEQxJjbr18W8dFK4RitR+lxMY2mEA+6+pZ6yvXM5V/c97XDw0C5ACsr6o/ntH0j1tq4PmHE9JRcxIOM1Ei9lBjqcB8wiHN6JgOChJjDGoRIEFEYx1KS1ngqMASywjtme4hKdeCR9PlD9RTqYRlawT+oFxfbbV2aiii5vF01ALhQAEKYH/0JQGQjGL1iqGEmCiGxgLg+FoS4BBbGLPrF7E/p9b7gowekXcTy42dztUXEdwsZelk4yAQXgGkqpoAJpCIRxBGhy7cTA4UCKhRivIpK42EXcj9wqOCUma2iDAksf1IZ5nATpFaad+52rgouoOd8pPCRmGYPqEZQdwOMPEYmtNSPzgwGkxod9wmjp2ll1q57n0HzPTyGKdDQ9xsXaPnMZk5gEfTb/Ufa42BdZnXl8vGImnjlfEZ4DkMEPJ4ivakf1iJWMIJYlSY7FEx7RYypBf1F3G1cHzPrOPk0cEYjcQITVQ8kB9wQMLCnC9z5wGZ7teLwbiHBtgr8RhIcRDMYUE3YfisIAi4MM6gJXnAWeITOiaTJNZAzyM7jYuxfS8yng9Y5XCPYH8nluJscBhrRbYArMbQh8VxihgccvmUDnM5AfcAysTPEGN413YHeHf0MTmw6odPauVx9q/35WeoEB2Lyfc/rgouAqNiQYYHDBfQ0FXIqHD70Dd6gENaw5jI2YufxwXTGB5uSKAFFfMDqCKwGJy3uB+oamODuKBabRkZrZPKDql09i7t1B8TGB5NBLCr8FIuCihsOUJYiz1K9T72gEkIKgiAmMgqgww8gKDZne8el+8Yn9LCfzwACFOCYVDGoQ2INJQBGc8UR79k+bYuzXOSBMqOZmfY/YVmboB8oz9iGI5GMYhTzHHgKxPmwEAzZGcjaAy3AVDeXRrEE3UkT4IR2rBCCCAAowqwUtuIXgP1ErRMjRDltCAeZB09sJhALXvBgg1YQRFZzj7bauyHQc4OpHFfYGfUvqAIBxfCrdQfoHeV5rZAEFurcwMsNMDENWIX/ADAJAbgw8I1zaEClqDS9mh1oXAJS3aH5jY7WiazoPrQ08wGDA5zxC5ip4OdI8X0tq6w6iQZMwljYSn6lQPgvnmSGQQ/KIl8zQBoBhaMsBRjarAawWaw8KeZmzBp7jeaXH+UywAD3gJOkJnVcHAHsRMJRXhSgq7j2+xcBzvouPnxEuWala4Ca+INrEL3ZL5rHbVMkKWEOFAvcXmBqoGKeaxMG1sLwDAPwEG+MxhFXLEE8IrH5Rpyxco/OloR2Q5TzLuPQA4WwCCgvWHJAvdMMoMeSvWH67fauR9k+RMokARjoshXNLSrljPpblEM5uIxbgDHvABAA19axV5zLUrLWHEKQNKN8bQSGqw8KoBxdyv6HAMlJGyYl0YBmNlWAsDHegYzGYiV/kdvtXBdvoyI6YoAHKrvQTSxfMRUMfA5G1fmqbRmhGUDKGEvQ34DykgClzn72gsqpEfYig5GKv+RKz8R40RZ8pU84XnF7jg+L4vg+iuTao8fSPpH0jx48bSPGjRo0aNGjRo0aNGjRoIQCqYSmkYAADer4gKNGjRo0IatOt0BP1Ki8DrQKFk51ChR4w5rqCqiJu+TK8a73YXaIULis9x7QIIQX634o/RCjeC5hhd4o0hcKgh6QiFKyxeGnEMBgKPGjRo0aNGjRtI0aNGjR9ICjaR9I0eexJ//aAAwDAQACAAMAAAAQkEgkkEkAEgAkkgAEkAAEkAkkoAAEkkgAAAAEAAAAkkkEEgAgkAAEgEAEEkAnfgEkkgkEAAAAAAkkAkAkkgkgEAkkggAkkEiWYkkEkAEkkgEAkkkkkkAEggkgAEgkkAAkkAE2gEEgkAEEggkgEkkkgAEkEkkEAgkEAgkkkkgEkEEEAAgkkEAAAkkgggkAAkAAEkkgAAkgAAAEkEhAAkkkEEggkEkAgAEEEkgkkkkkAEkkkAAEkgFoAkkkkkkggkkAAAAEAAAEEEkAAAkgkAAEgkAAkggkkEkgAkggAAAkAEkkAAkAAEAkkAAEkEAAgkEkkkkgAEgAkEAAAAEkkAgAAEAggAAEgkAggEkgkkkgAAkgAgAAAAAgAAAEgAEgAAAAAEgAAAkAkkkggAggAAAAAkAgkAkAAAAAAkAgAkkgEAEkkkkEAkEAAAAAkggEgkEEAgAEEggEgkggAAEkkkkgkkEgAgAgkkAkkAkEAEkEkgAAkkkkEAgEkEggEkgkggAAAAAkkAAAgEkkkkAkEkkkAAkggEkgAEgkEgkkgEggEEAAAkkkkEEEkkkAAkkkkgkgkIYgkkkgAEAAEkggAEkkksgEkkkggkkkkkkgMWYEkkAgEgkgAggAAEkgkEkAkkkgkggkkgEA5EggkkAAAAAAAkAEAhKAdAEEkkkkkggEgEEA0kkAAggEEEAAAAAkY5HZmQekkkkgEkggkgkgEEEgAEgggAAAAgEISoI9XvhYAgkEEkkEkEgAkEkgAAkkEAAAAEjgGsJ/3tSi0EkgAEgAAAEgggAkAEEksEggAA5YUfSrjc68gkkhkkgkEEAkkEkgEggkgkAkgjWcncv/AJYM/XZJJJJJJIJIBBAJAAABIJJIBBIrtS0P++0t6UlJJIJJJJIBJJAAAJAAIJJJABBkkUX+222OzrnIFJJJJJJABJIJABJJJJJJJJO+beu2DOW+0HagAJJJJJAJBJJJIBJJJJIIJJPd+P3tRkUyciCBBJJAABIAAJJJJIJJABBJJIFoYODpJWLSyBMMJBMJJABIAJJJJBJJBAIJAIBLhkYBIhIsWBfJJIBoIBIIAJJJJJAJJAJBNoGW1w/5INJJn7uVAhFFJIIIBJJJAJJJJAhoJJM01w+JIdIY/wArPIBQCASQAASSQACSSSQSCSCToGnQkCciEPr76JCQSCAAACSSSQAASSSQAbCQFD6v8AjyWazrySSSQQSAACCQQQQCCSCQICC6OgJIEFsC1eUfbSSSIAASAAACCASSUQQSSSAQT7NWemA7988fRCTLAACAASCCAASSCQALSSbSSMk9Yv4mk0t5JaTZIAAQACACASSCAIQCSCSbTJwi1Yhqbr3CSARACAASRSCQCSSCSSSSQCTCDBWk56tFx0XIaJZQAAIBCQQCQSSCSQCJYTAAaQTN96fPuSILDRIACQCCQQQSCKSSSAASKCKRMSTZfud9LAGrJZaAACAISJQgSSQTQACQYAYCAAAAnVUPPIBhKaQIAIAQQQQAASCCCQATCARZAAADvtYkuFLyFAIAIBQBAQSQCQSSCSACRiQAACCT+bskDJRZ6QKAAQRLAAACASBQSQASCCSSSSSRg7EKf25JzufhbCSICSQAAAQCDSSR5SZSQLaLiGSD7TL25UACKQSKAAQAAAAQbQSSIaSLJKQBk4ItHP6OIAAaaSSAAAYAACASCSQIACAAJKLbVs3FjQofpRCCTZAAADcAAAACQCIAIZBAhSJYZpjIb9B6S5QDQAQATTQCAACBRAbaSRQlIJDTgxayySZYSIBAACAJDSQCACSR4QLDAaSBgTG45dRS6C6GCySABr+aTgwCQSSCABJgKNbLAA3+0WctmTCjO3aZ++S23F6AQQyQITRJAQxJZb5arV/OySd54vCeyZgif3aDAAACSAbAABDaHTZMK6sSGjokk2g++bS6VBoAAAASQAAIJAbfX04CJdJIy4ged57QWThCUggSzAAAAACCAIBbdEZU05Sg/ujBA5vIBwACVxoWSSSG+IASBJSNuSEYGx6qOGdBRGXAQE2WAuECCESF7IAICBcbobbdzME+GXLBYMIAQdNrYVIAabQR/TUSQSbezeZ3YIDaalhCYbCAbYLJRhB72Dj18qC6zbcvmZNFQ3yg+QaIJbSRl6bBCKNjeJBMxZ8Xsyn7L6R/ViJLvQf9+TzozLgYmw0gccgASZQ7ugZZOWTT7T2Ftb2vbzTCcAiQbJsxDjJgFZ2ybBIhp+VH/wDkHqCkgVJO+CaiX7feLg5EfzjFwwIaZDCS74VKt4gqntoKAeS6T7X/AKcD1WcDoswDAdrZS08RxdhRfpMOkoIt+8kt3jMhchBJQ9gEpVJNd+V7nHG+tlg1t+/99vtv2ZbIinjPS4tnWtvd2E9xWCnxqVNXFlv02ks33kDhlUDNNkstowullEkT3SoUiQYIt99/+kk13/0lLn5+3AsmA0uk8X1yueTP2DKFk0vmlm20/wCtYKdtgsBgDamZPrUfPUGr9pQVbLzP/wD+6W7/AH9p0mV+Lunjspc3stnXXX5+ttYn6BVn329v/wB7McpIKpJ/cBCSQK0ZlUXnaf7pZqOp9Z/t9t9rLvhb7rd+ZMDkrfha5YBFEJ/tJpJLtvZ9Pt6T5Rht9/tiBsYDLNXu8K0Da/8A3fbW3f67T/bcG25cSbeyWUWCvzeXXBcC8aS76fzb/wD+3+232W8kt/8A7b7Jbh7f/wA5/h0n3pcf7abXf77b7b/fWf7f3e22z7Te/efW/S0K1pHf7+fbybf7X7b6XfXzf+/7W+67/f8AtfzRMNNui+2+3232+/8Av97NtfPtvp9P79/9/ZvCLqmJdsb9vP8A77bfbf7ab/bffb6/7bSbff8ARcKAP3dS+03++2322/8A/wDbf7Tfb7b/AH/2/n8tZYtgLF8qU2lvs3+323/2+/8A55t9pdp//wDbffZT0EzeAR4f7a2Tb/8A22/32O2//wBtpvrd9tpNnWnC8vEGDm9/pZtt9ttvt9z/APb/AGv2+239+/2/mAsJKw+Zc32023/++232/P8A/t9//Nv55Jf/AJQv3UYkIIt1bf8A/wD9ttPt/wDcf7/f/wD+n38s+2+xQR+AYFWTn+kmv322+/8Attpv/wDbbbff/fb7b6jS1sJIssylfbSfb/b/AG2++u3/AN/9v99/tv8Abu0cIki9MsyJ/a7/AG222++/2/8Avt9/9v8Ab77/AH05++czdhaNhu+32133/wBvv9pt/t9tt/8Ab/fb7pPf/cfU72Kl7/b/AP8Avt99v/vtt/8A7/77bbfffZD7/wCFxNSKOn++333+++//APot9tt9t/8Ab/ffanX79+sgiAj0Tff/AH23+3/2+m+//wD9vvt9t/vgdt/gyvFVhi2//tv/APb7fbfb7/bbb/bb/f7/AOt3+3Kh2P8AKhWd/ttvt9vv/wD/AH3/AP8Af/8A322322SP2/PPl0a5TZ/3+33/AP8A7fb6X9b9vf7/AH2+2zUO/wB6dzHSs8xdvt/t/wD77/8A2O22yK232++/+4QO/wBqpa1dmrk/s9v99ttvt/xt2b2lv2r+tt9X1M79Z0+7GyQlZZv/ACWbyX+i/8QAJxEAAwACAQQDAQEBAAMBAAAAAAERITEQIEFQUTBAYXFggXCQobH/2gAIAQMBAT8Q8hP8OuH/AIVcP/DX/wALon+HQ/8A1OT/ABOB/wCERfBQhCMohPPwSEUktlXCmXDHcaFE82kLuZUZZbw9mGaIkrhoSlo9hLwhvsNxkTWRwTy8Ez0a0LIjuKJZwJNNZHqSHrpm2W7iT3IbRVjAiVjZqoWBoxrt4m/LTPYbmEJXLGklnQ2kDbeWJYp3Hg7C4ahBMtCH+jNVjUY8qDUw/JoSrg32WhexDkY2RqODyjB8PZ2Fwx6gl3fDsRO/9GoRJBppx+TSiog0atlryMRahPsaGM7C0Lm4golTLYxyGquN6vJJWN+hGTHkMatAqQ0PA88djtx24XF7GCITMzVoSODyj88isRfZ2BJPpibaDXc2fnC9CTZHCMa6djZqBulXgTyMgkfke3BNngKyFpo/UbP0QtcKFawlCMPQ1DXFE5kjBJa418gt8OJNsSTjDMsbL7Fe3ANt9CVB8OF2Ma79Cb0Gib4yXkFsZFKIq5X3IuxkwVIrXUth/OWGfw/onNCTuviI/IrKEuDZsNSmBDGKhYy6Nn8GvJZIKmWQwhNnxpB+QfBQgwyvjY2GwEiujZ/OgxAmVxgwJrkZkx+QeOGXgYs3hkVNh9BY/Rv0DalHXrjBfwZtDeDefI/o1VG+Y2ThP0wiBMgmJtyuLZzOfspMyU2GN2H5Jo4xKnfIhP0Qhi2JtwxGo3cJSSNP0huvJ/DNE4MfvlJ4YkmsiBkzgzTJklonCFjDYUxSxRXs/pPQxKsfsbz5aOx0hi1oeJsJUzsy2MQmYkDbLN6lmgiGSJvLH5fQjTIUu4xMFrrhiMy+yCT0LcHf2FbmOBs9cPzH8MDErMBmTpjRPY+H/wC5ICmIU9IY1+eaO8E8Okyx+hDAIvGV6ilGy+fyUJMCJMhowGiFJIai1+z6n9h+C0JAWMUWjFC1IThf0F1XzTbXArsY2GYFRPApnTR8vy7jNTYaFlC4jQtoes/fgnmNIyVMUxo/pEOw/SI00Plxepczh+Dv0NYu4iUnogkG6Q1sbyiN3wXzCYjctkJf4Wmo2aQ9dEdTFyJxCEITzXeWh7/wuFZiBiQpRH/1cwf2cfba+EezGdcYpEwHYaJpm/8AvF6LxS+XZs2hLHCbg1Oy4bblMf6ednO7pk0v0eu4WHYM7r4I/Ko0URoxA38aI7BtEx9uFOp83r2UvROjfgdF5xYSfyh62f0Q3Q1SCpRI/Sh9E6dfEjZ28Ah80Qsl+SNkg8UZBLAY4Ym358M4nKGUfVOEPifdpvi9C4SGo9nYZ2GRbRjV0K0z8Ly+m8vpvVeE+b0T7U6Vlwx/4YewPRoYenQTadM2cU2PqvEJ8850X4b88ILhj4SoJZfo+HqhjXoeo40aLRMvx8r4EUfwTic3hfG/oa6H0LsWA6bDyRmgnBiFWmLc5aHEJ9DXFL4LXNLwhkbLPohzbbKUYMVSHgyLLf0aZov1l0whB9EINdd+N8ThcND/AKGfo4fGgYaDTS9jR6RIfv0F8VH0vhdF4vVBco0XidN4SrgsTYwKg0U0MQ9mYGYEyfXfknE5pOZz3HxSl4fwX4nxeUTUlhdyy+gtFSeRrOBtGofYwRJAEjT6aX4p1TonUurfXeucrnHK7YlQUgk4PIzJGCD0GegEnZ6Rgv4EQS4hrhfPTfOuUicX5KIx0QnGAvY38KNsSwKuDbo0SFhpiyUiRMtFwWR1UYvin0rzehl4vM5fKXN5RKfg1n74ySkyaCcgpbIRaYaf0uKXqS6L0X6i+N9D6mQWCOzH4NIrTwXJqehtBqccUFNQkbXWuF8u/k3wum8L4oTmcJsSpBafXEFRIzUpCGxrAnfojkQYYutE439CdS+subszGXoouJ3M3BcmKIaohUUP7xMj76J0r6752NcwhCfReIINm+GKhLJmUeMzajtbXZjOISpvpzh/G+f5zfkXTeKJWkJKPi99GRb4zQ8M6QlUxyH+CX+H1Ph83i9V4nyToXOeb07ILjZricoGHi5XkQ1sSjnFPRabF0xCKohF2GOLzPhnzXoYvnb6n0MwrEoKPCMQyJ5P2TQ40Q3UEtiVl7+K+AnO+O5rmmydOJ+mbP0PRjEP2KkLD4UWINYQ7VIbglko13C1XVei+B79OuL1wSG5RDUQmxb4ejQJDQyZTFiNCxvin0V0Mo/kXFGQgiC5SCHpsf8Ac52Hs0psuF0VUJ4ZtLISpMkj+1OicTrpgfTPi2B6SHwTtyhqITQ2Nx9jUVbgqL9E2Mkf218d+Tv1JGYtRFnlDKlIR++OBoCn+hUmxoTy/hmfnmFnsC0zsNW30Ma1Cox1skT7MILY8MZ+AUXO32p91KuCKx9j+s4k2Qe8pGhh2psSoLkExVsTASkmuDV6P+cx7ZPQ1HPLLULk+IXUJzyJ5kii4TYT0NVpDGOGoEyLYxVaXcVp0SOvLIeWNKJCXkdxPifohuK2X2VIglPYyamuDNQQ8GaCzyzBUI28EZOG4NUS8DEqOpBhs7jLwPSYuHauoc26E26p9+fRjB2tGDQ0jd9xtlgtlcJWJJbK64npFUQp0xeIWr+eVgoWKLmypuUtjafYh6Gp0Jwbosjyo2jYJMuHRvHzqTYeP7EAxJKQ3gQaHeE4uh0hThZQlZGhD/huXlUjP2PKB8B6GJlZQ3yuUJmYXchgsqFjISMvKSRCW/RNBqwGtI1dKHyhxsPWMhCSxI3k0qI2MWRuu8JtaE3chGpyhjFhROqORNncSMPmhRMH+eUmxMdvfvpTg3joPfGQhKmKSZsJHIIZhMH5NdjsEOqv9LYIWuD2dxL2JJaEgiEooxaaHlNFn8nIyqjA+uqLJY8DZqCyNHc0LYlF4EiRdxD3YlV5JK4JRGTMtOlDEltjTEjg9kzxsImrYhodFCXdM0GNZaGo55FYixeAvPShipvIhgPY9l4EWZJUUk1rHfEGglF9efaXYSbsfB76lsxCx4KxTYe+FqbC1CV+Ibl3B/0fsdvs4mxppIOl1BbGQs9xrORTuNd+E8DYhdx5T4iwesjQzf2J9nE9hiRjV26th5NhOxQ9lzx2C5Fy0fg9kDmhfsH0rjP0ZCEo4LWbKLdS2PKGi01HsfB6cCR0TIsYaFq0LXX3kX6PsHtxpvqQ2JqgsuCwuO9KN5vE2RRvE40zIuGvo3pvH//EACcRAAMAAgIBBQEAAgMBAAAAAAABERAhIDFBMEBQUWFxYIGQkaGx/9oACAECAQE/EPkF/g7wv8FuF/g0/wCX7z/grF/ldKVF/wAB/o1G5WPCNEICddiRi+bf6PxQ3ezSGq2Khr7KSOjG+zYN0tiVvQtiZOIV9/MtF2Nt7Y9HgQ1SaVGE09ISNtmyw8UJeBt8CH04NZ+RmnBKnsexN2E09r5boLsW+yrpCbQlWJzoSmkdDEeR4WGj7GL8GjLRPshPsvk2NFEm9sZ+KEJoTp0x4XR5HlDfhY3I9f6LRdh+r5Ojg9EU+jpaE6SMeEI84YxE3R7cOhC7K7H2bH8P5J4iJbGPSNAhQ4xreSz5x54IlVjRGiOxqqLR+/IvWdkKw238Jdi40qKLC4JJbYlekTSGxqvkexNDUB2gkx+YbIyEGoyszaE+D3oqDpyOsPv5B9Y7aQ3+yNNH9IM3QS4WGbs/3DQneEXbENRHZ2+Qa0IruiqIT6Kfwe3CTnFoO3+5fCUbRQmir8ZsvDTRp0jpNQmUGM9R8G1X6JP9+CdfBpDoTdwszK+JWMqR5SJ9EH0LoWONXcIi/Z1Z35vvGzY07WE1lfHJVcJeoaND6OhqjIHBtR0ZkMFf3jZ/sSMSujrPXx34QcEMJGU2LaFGw3Xh1Ca5pL6JSzojYvk7+PuGJUdGuG8XxuTayMaMPUw0U7v2xaUKODNsRtn4XE+Q6L6FaejqYaYVNGiCOD1A+hSiP5jL3oSrEkujoR2LlfhWLj0d5YVNbEdQQGN0JOsMYGqEJI+SYG5sgiGsSS6IQmJwuOi/GNJjJoZvfwfgA4l9iGNoaj9H9ipvwQj9FV2J2eKL0J8Q+Fw8bFNWAGgDGlUIY+q/MQcuhjX2xa19H89GF9Se4frpU0MGEhOpFGP/AOBqFH/tY1B9EOsrK4MXxF4PnpP9KMbu/MMs5q7HpF3+nPrgvYz1N+4c6pUKBB9iVGo9lD90eHyXzCPQS0xiQ+xyhI+MlyvOZfBfEJVZqeo7H2bvOx3ZJX56DJ6u/ilrCdIxLZdgqja0SLiEJiEzc0vwiz0d+ixth+F+jtl+yjEtzvoSidOr0eifAX0fPBl4IpTs1YSoim39zlMQUGUaNlzRYvorE9Sv2MF6MIQYsNY8QtQ/++Hg+7E6zeNV/nCjwyiy+c9LftLiEwuLGPhi7QkSY8hPYSSK9n/gxOEHwpeC9DrCwvZLk+F5M6ETS8AXTPIThrZ/5sTh17Tr2jxPQfG5fSSLt/wWI/MP2PudM8Mf/oO/Y34F4pcL0G2kPObUfYT2zs2/gXPfBcFnrMJzmGX3azeO48v1iRJYa2x6ZGjH3FhliHwYiixeV5QfsmLk+T4Ig9Z/QjcvLz5KYdgitH6fr4TDRSixeHWO/RmZ7lHeJlizZglR9cEIotkJpdlFfuHxmGIuKb+HaEQmEPMGibNv9sXZ9C3hdmpXyGkcJTK9C+tS+16LwpebR2Par6F/pYhN+RdhD2TGvJCftcHwnCewfqXDZfSeIM7PHF5JUgVwLRTsWmoM3EySf7Kj9z0XHnn16XfG+hvgjZfVuYTgtIG0/bFCTwdkOzFNJiqGJ/GGJnhluYI36qx1wuHxXo0voo6KL0U/6wSv9jCwuxbZC0dlGaKD8Fl4uaXis3ixZXCkw3m4uFnrLKd8GQQyly0NjVpCfgaG3oWF2LWEqho1gNU/BZZRjFmY3w3inWFzeELEETlSZfKcpjyNWCf/AFEJ/sx7ZG1o8C7YlY7NDVFov0pkMp2QmNZ7zRPjfTXBkOuN9DvhTvHWeoNghh9lmELXF3POAOv1DbXBHXo32CHz8Cy+L4LixcN1/Ro+xi0oeRp2EooJGzDFrtB25Gww8vC9t0IeVl83xvBnQ+PSGbbf2xPwMLbGi7EzsNVDwP8A7kKWlFj+MRCcrw8F9tPQZeaLzss7aTLH/MtJrZNaO2FMQtpBbY3o9R5RR4ft5i4vo9k9K8W6/Zo/oJW84RATqwhssLZFB/Qh0LDFzS+2g+S9CmuU9GChiZrySmLuDk2TJFRsCT/DQUVfXwUGU7z59K+juSX9kk0MQxPRdYSiaNdRLJ+ULJY+SfAX1Z6T0YyP1izf1lH9HklSNAhxEp+jz+l8BPSfPrN5OZBbn6LZaQ1OQtVGxDDaaHDoY+Oza+q/az3DWBOIJn7hitw+hMLSu2MGtir7Q0X0P4F+yo+VW/DWF5IKw8G6cH1lu4nGIcMQu+hUHQk+8PhPZ3i9Fn9cDM2GkPrD7N2Q01GiBm1oZQ8Pz3Vw+F9a+lRYmiN76ZYjvB4/pDTFijxSRHjEtS8P5iE/Z5PoZG+XlidItH0aLGiZOYLRSH4PIG+YC6ixmSMsX2QnB02vo64Wpom7ZoieB7RsL6ZBP1fMU+oKaHkWCy9HQSnaJI2yCcaPRu1GE6jIAk/9+XeMyiq8sQhid6K/oXo2d1SNtIfc7KOpDfrQzaDGJobCuvJO/tCKLyE6r8s8YehfR+Ci5o1dDb0N0GkKdJsv0iL2MSt19k0R+A3QdRAbWDKQgP5ZqiQmrD2OdlFKfQkhNWwgX0QgTPsj7Ei6QpJI6jOmjZrZqxZPz5Z02f0dCN+Ma+wkEvhGolQTK0Sw3hHeOzRXTDE02LfYavlR9F2EdsST8icJEQmJw9DFBsw2wtyY6mh1hoy+17nXvKbG02hu40vCLwJNFFiZgxB0yQNENlDuRH9Pc795D9hK/wAjIvA17C0hPCxN8HMaNAwm6S36SYdi9vfeNFfQnY0dl2xUQQJObQ0alaRiXZRY+jGi/k2XR0EoMfmhMuxI/RYrTlJbOjGH+UQajH1/R7afsSimGqOehMLlieG9j2oykkWrY9WGg8X2X78nUEqSEkvri1RdlwxFETaZYb0dR6olR4H0fJ2g8j5grsZYZ2GLGjKY9aG0PUZoIbQkdIJ+/J1dfRowh+3Fi7JRQ9D0I8HnDWB9sTjQRdMk0UAvYT4FoqUbZrHIxiDPpCY3RdY84tMkO2KKR1IWXYdpJjVX5Ggx7Ei+RKcXgzS0abHIIXR9ng2dC02mLoJ7kuxsZZfItJG0kTFKf1yfQuzsiOgjwPsbwEoGiYcyJtZA+R1wmmbZvHJlCNvvQnVrDwXR5H0zpZd0aMzjwMee4Vxfs2Pf6CoYlf3yZoK5o0QzweDyeGdDGoJJQW0W/gaM6/2veXhv2FljcU6lz4Z3fAusvB2Q3UXQ1RkgjvWMk7PkvtmsTPR3xS5Ti0kXRYUSmZli0NOVG4qNnjHYS0USYgSbg6hIaKaCTTZC+/R6xONxSlLj/8QAKBABAAICAgEDBAIDAQAAAAAAAQARITEQQVEgYXGBkaHwscEw0eHx/9oACAEBAAE/ENMNweBzCLl8M7/wuIt8Zeh3xv1KzLjvlfEHMWovDKLcqlKDW6PeDcYZcclsW+O4OeWGvUej9R49A9cdQl5ly79N8Bi48JfAUcPpa4Nc1mL4mr5dxl8JcSphMGF5jPeZeZ3Kk66gqGYTU79ZxqHqZ+g8QLlSswK9QVy4m+bjXqqHCXKolfWbx6Li55ccVnkx1G0oZaJojXES4KEIquCD6AuVl4pJmMueUzftFqDcWLP2HiYY4y7/AMTOoN+ms+q4N816Ryt8kK4DEMwxd6gK5QxIKihEOHhZwA8lxb51BjmB9oscz9h4h/hxfC8xmJcWGvU35alwb5q4uFudS8x16DMqiHJZCSkGozSNRa5RuagwQlxai+JfNxzKxwmeP2HiE16rrgx8Rm2XbHc3wNQb5VHDLjliDdw1NPQvBxol55C+EkMQZv34vHNpHUdRFblcGOuTUvmpqXLgy8S4tx9p+w8Q9S0RhuLl1DPA2yoPKlxebxBuDN+hqMritk1KuUweODmUyrgVwN+hQ08yh1iBYG25lAm3iv8AFqdz9h4l1qD6V9TwsHoupeN8KVDMIYNTAr0YT0qzAgXArhPHN54NcsXE1As8y/qFYVlQHhUly4N+q+f2Hjg3XoTONzq5XBzrh9CoNxwS4uYPBSTF6l54WoueF64Y7hl/xHLnhilyhiTB3EanUu+Kblwf8H7DxwNPHwiOOuNzXpq/U6lU8jcGoo8nLKz6HUIedcLRL4quVxLxw4moMuYShlcJEzAiZ4KfTXP7DxzcYSrm+Wupv/Gzcqsw9d11D0nFy8cBX+B3yLLvg4S5XLA/wP8AQ6lY3GENmGpcGMuVj13wESuGDEoiVHJBrka4G+Lhn/BtFqLZZLg3zceNmJ3wPnjvmqmv8FxyntP+EebIP+IxwwYHCQ4040jHqH4ilzfDqK8HFR4WiWj88LqXwM0l3HHLqDwb46m5dTcfWsu+P2HiXfL7TTm4s/KD6GpXBcL6TmJc90qokD0h4XftL3FXEcsqPFMqFPGSXPZ6gjL5WpcSHKzIl3Dj9h4l1wtxcIvnTB71MIS5dy6hDcdR47l8LmuK9KZiRjXnjXO+L4cMLhqJZEInqNc3FWOZqEHCqXfp/YeI7l1GddwgvyMuGYsGMSBwImJVym+Ne0q+DLK4CJNc7iYiYhr0a4sm5XvO54i2S/VUM8LUuDyOZdnCXKzD0fsPEawi7iZnDJuGZETxK479B7kOKl5mY8KjiDcPQ6jr0MfblYZ579BJdems8HDi5d8uIN8+3KU+j9h4lV1E50ipbEb1Cu+GmZ9JMidS+N1HEvURua3KtjCGGXUG+HU36G+d8PXFXK8T6wyxyRfM79Y8dOV8MuDxXoS5fP7DxG4SoYgCA8Qy16Ak1xUC+azx1FxxUr01BqLHJAolnOn25n5VCNdwmfuU/MLI7xJ+mUoHm348EXrphsn1nLO8hBQBu2P2T+YywqAR9g/iFAGv6Jw39IHUrEsYYJpH/DXC16O4MvhxC+AvqJTO5+w8R7zMFRwwSjhLiVwGYEWsQyemuKhj198MXxGC9Sv8WPyRHFsVWdY0fgZsAcoB9RPsIpF3r5UsqTwQjKAJerFwttdQm4HGYvkLgCtM1yHBWIVeCi0jrZ5lfLFCBFadu9wkXd6BCLoVrrShq/mT87IKZykKEuzIq0QRwswZ5VU/RPiUSjss+HyfxNw4eBud8WTfcWo8N5g+8G+GDU3w73NEXxBJ+w8Q9ksOApgjyl36GpdRxLzLh/hVORFhx/zQV4Nr2IwkJQ9eK1fBnO4gto4KgNu+O7fYl4Ad5bAkvBsLZnqVt/Fwq6p17PMx8pmwOnhWwOYnmgweCgAiHudmYbYeRdzwx+Y247E4MXKGiQ4dgXgaTAN/dp9eZaNn3R3TbbOw3GqVO4ocVS3RnbcFjBwUO5vdm8udyjyBuMUDFgFbYdUw0ur4DeHrzsxmo6FjKHqvX2PaHBIQW0iYYOYr1Bg5bQKImJ1ykZdQeBlrUX2l3XBP2HiajuJcMoUeX0VXoYdS4bS7g+haitQahqLUSFSorvL4e1+kN3F8bXkrA29uWGuyjlKFPh8fyZjcbZFCLr22L3DiE+vsSYUmrXtWGhjYhQQFJYjVJdykBZKwCdK84qP7LRag8C2vpCnrSgD6RC04Xc/W5XAERAs13BJIKHPtNy6kIpku8f6S0uGrl6migLdDqX+WtozttQ6yLFvcCamLF20Hvai5l7wlW3jJPJeU0MsVi1XntKt2W/p5q5tZrb5ZFvYy/MtvSH5A+hwkKaZXpqyHj0FoxVQYalcPo/YeJeOcsy8pXDwlx9GpaQxDMuDBrnCLBiFktvP4zcv0i32KmrFjR4D3Jg/SJpZA5v2EuBxQ6nAHvUcKcio/NbWDfHxLvflJX1lUFDSvTW6+8XGlrtfrEMAYWct+Cd1zPJXtCDvVfJXUSYA2XbTFH8/eO7SLas1j8wwQgW4bUrsbz8ysUoLoLdH4YASCOHFjZiOyGgeB4Tr+PJGG1A7/AA2y1HJuo9LqoDDDLOz9ItRD5kbflG3rm3tdMWAx7Qi9U19D7DFMHfkHQcJ6bl9TvnfDmJcwmj0XmXjEcJ+08HIMCVHDwwb43w6iUTccPF54uoNyoGJlhElEM0jky/ulaD5lANgC2sAXgN+WUNktunFjI7/6M0Vn4t6n3ayUw0Qr2oKzaxnVUb+DCbMAbFBgM6CUrq0qsfhltsHqWWtvlzKFXQqpiorbW8xfuMw+iAUPeO55Zgb5fmUFQYoaVrE695YMXcT59mADxFZBblVhjxvJphQud8F9q9CaNzKvNaVs3WqbFVc31KlhrmLgHhYPoeoLYFiWJ59FSv8ABVxKg3y7juDU/aeDkGHDmLUc8XKrllsMzTPPDCGuHLU1xcZLRPBRm/bU97gbL0AxIjQsIfY9yv8AE6H0MnXaAY8Q/XBObMnr2Ya8bBZQEW12yhXOQOyCQeN9pUp04m16Rm3w5mQfFTr8wfqVDCvggXRGysXxMvrC1N3rxPmKtVda9rCjjYYD/wBOnqNja1B56mzz4+kp9VXnwsQ2VTbwNYjwzhlGxMq0Gy+zwmP1210/rYLe578LUWoNxa4XPNReuL4qJDUYlysT954JVRg1B4XmPF59pd6xL5W+XKRs5IPDxWIkwQt8cffPwMf1qRbhPfB9l8Qkdoic+K31SzBDkoHeIACrgcoWria+DgDoVoAAiZwvk3/uRlNwti+YlXXyShxpyM6eWGbHs1HPxYP5Q/lL+5hgfLiGM+P5gW194teDAS8EDz2DxL1Cjt0Su44KrGzFhe6zVwlJ04pkSdhecU9QsyijPbshJT7PuiZmMIC2s+B+kLF7i5l3Bg3xXorio8JfFbghP2ng9A1wG/Q45GLv1dwUJeZdxbgyszIekz0bvvPQWy/DuDJqMI7HGhTVRlo0c2kat1xAhC/9CGIawAZxe+mfRQPMAbHLUWt9PzBsy+Jsj3DKlbIoaNzBru5R1ESsT2Jg0dfmax955fYgKc/LLtadO2WOClpv6IM8bXEFe0Bm9ppt9DV7IGg+Ljk0htfFC0yO1wEwRBu0U+uX1mblQmb/AMV1Lbi28LFpg/e6PRV83BrhLicV69R1KH0OJ7CWqCCDUiRIEUA2GSZWB9Il+6yi0fUhMRkwuug1R4jUdalJB2V5u5a0THYxoWWfxK3N+CZ04S5hcWcFT3o2+xRlscb6ytDTFN795oty+JS5fuxcUGJR9eQiwC+1cETEL4rbiKyqAvO5lzOqyFpJQfdEsB7Q6AdAIzvEC6MOTVcrUvhYWi4l64ZYn8zuVm4uY2n6Z0f4Ki4c49CXFhaM0R4WpcvhhYqwCpdY3omCzG1KotaBkjLqKWrOxaQ/qfJtI/QxXhjStMp4nymBRZ+SBHO7/cwQqDcTdx49GvhSq8DK0Cr+3xEjVWnmDkZJly6l1r7w8mj8xGQD0bYutEcasO2m/E7qwcEKyFl/YS8ClEEuIB28RExfysZU0h78XUeBjU1LeNdyrnfFUb4SfsPHL/gbiZ5b41BuYly5c+MQxLSPxCYZFGEtDyhDkVTIvzBBVyTGqU6erlotDh0Zd0vedhT4Y0ULPeF1taZUg63W7/4gVyXxP3oCEEUC8/ccQU5aJfg+srtx8y7f1GBwd6rLBHfUzTO83bBdU6ja77TgUWt1ZfmItIKtYUr+D8wKl59uHPGtxanvN8srm4vAz9h49Jji4tc3Wp3y5IQtPovPpZkeBdyg/mv2iI3l3VGS3RvqMPfRvUUeUGHs5evvFOh8jMb+V95glUXoliFVUq1beExja+0VAp+wvFb4JjKU+Uf3CE+x+ryFgNrUUFtLRg+iYOUPzBFhb7w3tOj4vB6hfSUUwFCYxj2qETTarqRS7eapzKIJkNgf25bwqTTGjLvJN/PG/StRzFog3CXRP2ng9fdy5fNQK5biWeJaa65PTXarfS7D7/hQU27RiJzQKjZpjGK1EQxZDkuHWRNDGpXht8kR2foz3JNvZAbFa3VH+EYPyQezn++HcDMFowmfFydR0z7L/cHPAiWBf01+Zn+UU8SjuT3fYljsvvElNKxcBjnN2+wwFYnugFhCYNdoye3onWlySBhgXu/+Ij6cmNvovhxL4XH1ftPB6bzGkuLkl836KlDAiXNrlEcc0+Jk5mTLFBdL0Pl/YSrWmTq26BXCKN3KpFWNzYUALXXxLAZxURQcd211ZExOXzPKvvUVN0faCl3iJJkDF1a/1NZoO97J/Ub47nnwH7/8ygfGfB/uBjhW7DVX1f6hUhwnyl/3FP8A1Pk+8ASrvzGgJdZxReWxoN1BVzhRUBFloMx1iwjDLPa9HuIbkM+gKD7cisCvUzfF8MOT7z9p4OWLcuLCa94Mdw+8yWHoqYiVK9o7juWlY5aeYawOEYa2slZaj5xfaCG45HQhfc5DGzJNgefSonAjfdhlqOQYa3HzMyWKjwStbZV/S5cWSwL8i/xPBmV5p/6jqPUvMQHC2Pd/0mjhSxzYjrL5NH4CUw9qdXj8T3F/Se4S43wrkUHmSgfMBKHh/C0KcjjNkxAFmKbRqhtpq32lepx4DY/Xn4D/ABLTFs4IPqI/YeIe8u2ovXFS7lcsIYgVw49C7lxfeU3LlXPbi4JliLRjlfBXs0zf5rRKw8q/kveJdSTs7x1C83nt4h6dVjX2D321juIdr4E8C+uYWtAvZt/czJRI96YIlsZ+FH8sdR6Ib+kVLu83idvvDEgcUBHatENuAhnbSfwjadm2WMq/hh1RWrGo6ANQBLaUzcAvF5NR7sIG4s0SzQNPGNQkWdPleTtfxbBvKNoAoA8BHf8AgXPF4rjXGvQQKn7DxNwyeIkuuO4PpHcHHFzcGvRRwBDDFHgV4ABZZIWjxN+Q8xjyiB/G117d2aBGhP4LRg3VLZeWqItrSKLK6f3pg4MD2itQo101AslVq8j/AEMQNl34SAqkp94tTN3c+bh8Un9xL95fcmiRKy0vsf8AQigqlt3m/wDD7w6D/cOhv2YbdKFhl7rNPdZ67uLPwAGYtQ4Hu8OBwsvgYehxZ0GaO2ZpqGzvul+2pkm4ai16biy5eZU1N+iuX7DxwO/Tv00XD5i3Bl8DiOUyhrj44rjUS+LkxnUbnwrvt1Cga/rQ0oOnYnZZHdLknTbawBbXXm4qAxdHFpmvNWX0krOAvARP4JhREbsaz+IZajeV5YNNgvzNqzNmszLXZfb/ALlGfkY+J/UQEwSstZJ27a+n5QF+Ln1BhihkO1MXD8M3BhZYjZvDUbPlHCU7/wBFbbomTgCEXl9jQywoqgAPIT+DQQ3EuVUNem83O47mvRUd8VNEDj9h4lZ57xD0pfCXGAw43DkczavTd98riULpm2/gu/Zn5hNhZF+VpGNPjUfZG1oCFTIGhVAQGqtKytnsq36wCUsnWH81wDxQT9DqADsbfedU2aYM3qjwq/3DkPygqfxDm3eEgWtmBih/Q/eILSiIGD6ofWZlMhEYX8giRFISZKcbdtpdHa7uNWdDCGwFq+WfBAjjVJb2m09rKt9L7Ssxvga5v0GZUC4bjz+w8eivVVf4xIJwtRe4Obl5ipeJqXcJT+HHyeH3My5TOHJ7bj7vmNtmxiLcF9juLnQFQIHzLRaIlrq0KLiy7qKeMGStYUp0vW47RO2YdQd72Ff8sJQda7NkMCTTH6bVXzHEDpCsgcvvLINkFCxBlunqdquVR7P9ETTyqKf2fnl94UEMvvxT0VmdsWYlT+Oa4CGpVTUCuLxOp+w8Ral5lvmDFUXJmd+pcQZcvioEuiaS8Xxmdc1yEYIUlwrmEU4IUeuFR8ZhAblhXHuRAYNCZaoszmO2vxNj8RWO2V8D+oh6zBmlNERVx0yLA2D5C4l2QpTzNVV2lYJVTL5eX1ZX2m5VzXBk4q3lYyuajqBngeNRYuIEeP2ngmGXKxK94FwK+PTT6lwallwb41Pdg3Kp8x3Nysz29KYY5miSvaB/BCNRaK0iqS4cw1YQ8W68Fi5irUQJXzNhC9+/1Ux5Dp+TuHlBBjtrX+ogvpJgrMeMMGp1N1wRhri48M1K9/VbDcvcufxFl3L4/eeCXyemuLYwjqd+m+iDDJBual53caIzuJngnfDqFdDXg3rx8/eYAhwPBVEaOtbXYgFddt2yilXGtx4onYV/nf8AUsmiop8wvmK7zLkIbJOn/am5shiXZA4MEXhbgxmP8Bw41Lm+A4/aeCPHf+N4eGVLonW4FRwc3xdy4zqKQK4HG9N1pP6WaTBWyBuiwl7azMG5sr9oinNqB1BbX5FwwWi/GJaXZ7xR/iuNw3LuWTvhgSsS+H1hiBcWuAvi4ZjH0v8AwOHWoNHA8am1l1Bt9DeYXHhLhEuFwb5CJfFYlMriuT/UEYrN0UKyqj2yu4HairdYG4tnP0ju+ujUe06kKnqZZtZCqJhyHHeMSi8aH0cjcOFqLfczOpcuHC+nLmokcPGpWOP2HiVxXHcGuCxYTfoolJUdQeDUNf5dSukfzBkswL3AWFnKdZN4gOsxtzSupVKyYH1lf0gr6Jc7wSiHNvjph2aDFYRrTPYA/gg1CEumWy+NxJ7yp3LmIalZmTCB6Gbl0xPaDTMM/aeDhmuLm5XOoNQb9SQMymHj0LXoWD6NTOr2/kgpdI79mIosdS7AdKLHiVS7zBqxfb8xiGmSKw6QYEFbs7+YDLEC3Sv3EVvyn4mupc11DcZWY3AZn00QJUTl51HHx6f2ng9Nc3NyoZgf4CV6e4t8XUIXfGpeLh39WfyRO4JTBKEa+sAGgh2/6gihj6IGu8v8sPDcAWNDFaMQYlGxvLz7QeKql8NQLq7e/ojxdxpLuXDKLiGuF9Bn/AxfReZ+08HpOHgKnc2+o31Ai0S5mF98LXFXKIlSreLZb4jLmXUAiJga4mfMZ6UFHSQPzHGipTevuQkwf+EXBaKnGnMctmWggtjcd6rS+p4NSveazKJ5niXwG5WeS4a5tl5lykpy7hmOIxP7miVX+E3UquCXF+8NQi1NyoPG2JfDfiVVRfaVcTEMHNQHaDuqDDMPaTMfNgnFSucedzR5fEauyD8JgaKgfxEEBSAgW4PIedSz8oO6eXmZ/uYSvHFSrlMrKOKxUVdQb50zuXMJuVL9KXAqJbx+08HIeowlVmXUX7QWLFhvjbPpCuAqXPiai1FzHXCxYLlMjqw8dwdUfykvnlk9pAIWnn5dZfRVVn6SqgkBKwkygBW3ZodfSJXd/wBSVqVwN1AuO57RKhg1wMc1xUrN8p3N+lhx+08HNVK4VMESZqXUvMXjTO+L6huXXrMDPC1Ny5cdRYBA26N7JdP9vaXa7yvw/wBJVmGLP7LKxvIfxGptYf0hB+WRX8D+ENQKvjthExKbjngsJdxuXPni4+HC2LcGtRyXBxLuXiXFmqn6zwSq5JfqO4tvFcVUojmEup1D7egeuLi8bcupdW/TEweSF8o/tBRILMFi1uxt8xcYlisJ/CZvd3ijSVKqq/jzFlZFFT6RH2gsGXFhqFQnmEZpiM0xYtkvjt9GpcMS5UZ1P3ngmoQxL4tmFwVeFUupcIz35NyuB4I5l3Fp94Zzyu2dysPDMnV/sTKAUXoAtX2qcARJDQBVXbPcWq2ZUFiWqsddyyWX74Q/iQz8vTfcTfrqu/rFv4Vu8SIb4PzO+EIsPMZUvhmZvjXPcOp3w7uDUvM+Z+08EslVNseBSOWDUuo5Z9Yw1wMXBOoZWHHxng5dwcRmGMMw1w5YK7Vn2IZ22+/CfkQ2HvELwRVkLi8dSobFj5v/AHQrlJsopFJY/WeJb7NL1m/7hCEGmOZqbnfFy5vjNf4DMuH5jmdxx/uM/XeCWhn0hXFSpXAeu5eYS4RhNsdYnUWJcDM1wu41fsH1ailtUh7K/wAsNd/SLfseIqFtWx11EHSi+hf1GC4CnnEHR4mYSSqAa9z/AKeCVCBXDPpMw7h8cXH4ie0q9cVA52e8qdT3niVPpP13g4WouZdMH1XxfoSu4Ra5OLvjU3mdRYNy6hmNw3+hYkPQv4P0h+Gqiwx7s6ty5XcwUQopoLItVeWNar2711BwidWa/wBFKktYf0/9lovhv4gDVd57I/1OveBUzNUcBvllRaiwg36EqagXKqY1PMvhmyDc/XeCDGXUcwly5cYvM6g0suXL4YZlHpN1G4O+H4RhPeDmXDetafeXij2Av/hLl8bSraiGgMtqi6pPNJNcur1GdLNdcZusbuOjt27NRUbP0KQX9BIXl58fMbvcQucpAwyfNoifwzxxrgIFcpcbubcEDhwQb4dy8S5cZmbczNag1LufrvBFh8zDFqPNRuXmV7yuRzHftzcWorOW7iy4xl54rgLJQTZj8Rm1X0xlp/Nwpu7KYijhTae491ssG1bZYhpAG/vHiI32Rp6Z8pUKHzVGrbArrtguhmKpFWHn+DNepuXVE33shrjcITPLKzNpUwS+dx73wZjiZh8w47nfH67wSszFT4574uXFxCWkGzjXcG5hLg3Hh3qOSNJds74XjMzwNQCoo26if2DFWIvYq+ks35Q3sAEfbOpVC+CIE+8T9Px7y++WOmG6unRuYDaSAdI1nzUMW4ZpMqaybioCZ3pBG7iEDI5JuViVmfzytRcTxKqXnip3ww2nvKmZdbmJ4EW+pfBP13glx4NxzLl+8vi/efMYZlVrnffAz4ldzW4sZrjHFyoTdy4iwOaCq2v4qNn8WAUawOi8wyYlhxv3iNt7mjX6WXa6fyQf2gHQ1pcrVj6sUGvYi8d5uMgjjNju47Kq5e7Rf5mYJU1Ll28LmXXC65B4XHhmiXqOZgly8y4y4f1uidcnzDBNvO/QYY3E4GuO4eEvEd743Opc3xVegNCZZshU+lqEacvo9Hx+eUeZjLektTSvfUsf9zwZ+YWjQivvLkoUPmggLDjY1AXACHlJ/JDbQ03tg/lTEPHHVKvwkCMu4/MvDPfi/GJo4u48XnM3KzyUZ3C53DUsZhC0W4u//wAiXTL9B9pXiZuOoPI08XGdVKuBAZc/E7jKb3KmJi+Al8CDLMj1efxFOLPsUKhtZZ8Bn8oqkICoV3dX2N5WozcsVqe6daG/ue0MUYjdjZ9GoCS6IpDQznx/7IzObHiYEDYrdjF2bRYK7S/knxePwH9jxVXNc6IPFcXL48INMXNzfD5m5cWC1Ll0QZ3P13g5J3OpozAIn34Ri8jiZZ3CG46l4hHccVO5mXmXbwMvm8bV2fBL5aFL6L+FywxQB5zfzFEmfiiVsy0LGvtGYhhD/QLgEVCKKT2gvRcUKlzwED/MMGzTX0l1l7Cwsov3QDmg2UlZ7JB97VweFrkNxZaLBeKlehpLYt8O+BllwdS5+u8E7mmXwQg5fEsn1jmYSUeZUHHF5hLOp0i3L1FzFg3LwTE7xDU1CZl1O0sJ8v8A2fRR9MH8h+kEWiB4CJZPZFZF2hMtbZ1cAu6vSBsA4S/MRzaoB+hiCDWfaV61mPgv9Q9gGGMIsDs/LyEy7xA4JqifD/pzFScJ/W0ELxvES4ko8xhg40QZcu+LqOUWbI5OPni8yrnfH7bwT6zxLtl8XiGSZlVDipXiBKl9wZ3LxuD7xbJcvhrfBklZ4zHFSgViuHCA9pfebm6o/wA3ghRQlmRHpkaNr7JfEguAvV5XDo6jZGMOodRCEOiJcdZlGi5Xu39zJqS1ow7prZ4lKiVCpcWddPCRVm1BqqAX+IIal54uJcCJGJL43iajiPFQudxEhKvi4y5+28HHUPM3NTE6jDMKqG5XfUaZU6qY+nFx1xcs4GUeHEuXL4ufFKaLgl7X/wCRGsqftYPx9yOCBLApc1KrWufLFsIjOBA/ciuu4Nq/MCY6E/ojrDEq1OlbAqfaNpaKjFWt5XwQw2cC8XzV3lHV0P4IfRH9xLrEvisyp2xS4tscTThdy5ZfBKqDKhKpgcMTHiM/S0TU6iYlzRDUFnWo8WwepWIxmuVWaYsPeBzdS4RxFvhwagmfEdOiNoev5SXAIhHug/kMJkAFq9R6y7yFoN5UW5BQXMgtNQJo+MF95l1RKZgaw9kuoVwZ+hLh2mHM6q4cvoJhKokCAv0v8zAmQnxbACM/QgH+2WPQX+z+uLl6l541FuXG7l3Hcv7y88ldwPRVyuKu5VSmfsvBxdS88BBzK4Uh5jmbjA4XhMTVSsRJWJaysRzO53PmO+HzK+rpNAB/5FVzK/VpQKulr8pb+VhIAhSJdkJMa0apgwfHtLGdH2meWVxZLgWaP4ItQNRlSPj3BF0R/KJWIYPL/wAIe4bOE5xeoOaFYTGB+IZfJcuOY1Fi+vOoPpb8RIR3H+t0cX7YgXxe4MWX9IPncX7cXWZd8HKPvxc2wHiqnUdT45I8M1iQCylp/EUSOcEQUFoK6wwFAUEw1aJaFrRnREphTMvni0Xk3EDdMggBLYXRbhuYYWjoc7JUWW2G/glgp3Co1faeIzqg9ZYY3gVb4gR2aeSj+4EwLmzajH4Z20YPfJ/CXgjnio4jGPH0gXwSpVwMSpeIHBNTUvjrj9t4Jc/ahdQyZ4qmbZiXjjuaZcIypqYZrgzDLHDGWS7rjfFXDT0zAI9QdhLzVNvjP9OoRjhQlK3iCqLuBhlz95m9YO4W7q9woLc9xSP7wVwxHwb/AAjjd/YwE4StXmsypQ1Lwqv5IDMlpXuI/wBvBNdRySpt4PARKlSpqfEuVc3NEM8XmaZZFvj9t4IuDeuCT8TUvPF3wOJfiDFl44N8XmGINcLK9pU3CbJmFTCSt1eZVqLdo01a/mLnKzT0lPtFT2PY2KKyOU1AkZJUKFNWNpkDasx8TmjbRYD7mcwZrCNMIMW/PzLSo73NHv2Eud4pCqluCihcKc5DkcuEgEQ0NAC8/JFrbV3yD+a4GtwajA/WXiOeDbBHMqo7jFph8QJ3HEGX95fJLn7bwTUNQ1DUZQRlS5UxxcJ3xVypi5Ve8vEoZd8VK3PaaIkYvDP0EZgFrX9BSAUMtNdafjgYba6LcJMERYmpdMC1ouoXemvMv7Kv3iaCV5v5lm1Y7jImpVLZx7zR9JgWL1YfY2TIIRM4DJKEe3g/nr6c+0r0tzj4DDIeIb4vhb9G5cc8OI6jogyubl37c0y6n7LwQG5TDUGE6iS73xfU1LHE75vjR5laiYg3PedYmZp4MxZc8x6iVSez/wCygy0B5F/kQY+bd8oFwzFK1qi1QPK/E0JE8wwZGl0HzH4Slk1tPlAFWxvqFAbA/aZt2+/yywnpInK3yGaWrVWeFS0azSQoPFs4689abPadTB58UE7ouzx1G8TLJRHPwQyGz7oS8wqXPHC8EfQsuzm5uXd1wEovccE0StT9t4Ja+ExLlYuEe+GVHgczePReY1U6lTb7T24qVLpjGoCLogMNkfc7gh17qd7+T7wVwxN0o2qgB7xZhVMQUaYFvRdeYc1rHDXmF5Npa+ZdBvK/zEp+O4/0agUzilOJhypK+/8AUNf3BHBPF1ABcEUV00/7nm6x9ES7jye01wtQJeeF05iy5cGLBSXwLMxLl9QzAfvaJ1cZd8XXNzbw8BUvMvnxLxDMqLWpcW2eyXLl/eXMn0DzOvjaMdkWh4ofzZFItzIfIgFQ5dDhlljXNO1VTpTS2XnMqwp1aQ5buxjj5qAIzBtkqt/d+0DfPf8AcwQliR0xv8hoW7sbjdpgPlp2If7iaJQ/n+pZlgAfI/pGN6ob+RlhVPVnSD/uYRcy7jh9Fy6JcvjMXrl4uFyjjUvMWo+z/wAiXibmhnUubcFOXgyQWXOpcupdsLRCS5cuoMuyX4i1BIDN71eJsrX0Bb/DAtAc9u3+ZGX7yxyjynUuwtjGZWQz1Etk6ur+sBdjZpFUOhFEMMa+LsUxLmwr3U0PaJIDP7aqOnUeCWkuVR/uXQJcKZHA/mE9kq/lEzdBfA3kf6YQAoJ8ij/JL4upv4lYnWJZcWpcvNTUdy9xcQnc7lalQLj7y+p1LzmLP2XgnUuLLzxUuoPC5fDBi4l1GbzCCkGpc0iz2Mvi51PFy/YiEIwhvEq+izo9R/VZ+K4uBHgCayq1hZhTWASikAFEBySzUoEsbpF2HCnmJUAAMlgf5nsy8DhrEMmRLwQYuWG5wVBIPm2iRTVhleo4pUr6PB7VHJ8zJlfR9pXxLe4+50D+Ge86gS5eZ1Lzxct4YxhxWZRUJdnowyvM/ZeCXLiy+5ctl3wnNy8S/MFqDFlnUYtl4mkuOXLB64DeJdYl2TJJAC+f/SEwKL7Ch9z9oTmE17FTXF2g6RIcbJhSmI5oBbsQr2xAOdWjOKAQTuVdsPhWHKLClvRDdaqvYGhuqW0dqjLqOovOBtmU/qriBhyGvZDoxkMVo/EULiVayCe2AxJjwvYGTrcGQBk68n3hDXnm+Fl8G5cZ9Ybl80xxL4Zc1mYPifsvBHCLLjD0pKxL7hUvgfvFIzcvxLlxl59p7wuVTAnSNjccHHXuFWDvRiFVCYDR7joRmIO1omVJqKz4TE7+fAfxcIAPPECuwsGquOz/ABVsooJeTAwYyWVXIHZV1iFK2oG4UKFL5mrjkDRqrPruVYm24ALMmDNh8xPSED7pGiwpi3W5oT8dQIFuMRDEt6xsw+AbA15ggnayLE18BGICcQCLRdGnUVBoXxv0XLuGppncYNPFy8wZdwbm5qdxZcufsvBLl3BxHLLgxeFoiy0u5cHi47ly7muLiwhAuMJXzeiANgLVfvtEZSsbGUP4f3h5sagoPHyn2goXQpT28QwqfwhVkfrvQqs4xeMvU0l+WgfBQ+0u5KyZD5F/mastZan73LW629pWvgSX4h0HswPqww8ZEXGrD3UajSjmUzKyByv6lng5stp95Zq9ojZ1am92FMdS4MdcpHhiBGhl0wblHmYIVBpix6hHyRquP2XgnhBvDHHAYmoRpFuLHgJqMr78aize4sWoblDDBAuBGoC+Fo78fxG3sUa31/UBSrYL1/1jqIgJvd2Ms4NKIX/cqAJm7r7sGkFaT91AEDW/3yQkPYDv1CvzESbpk+1oGdLSX6qH4lUY7ofxH8xK/f8AoGWg6NzuAaQtopcySHFCV/DspgmIG0fw/DUoXCsHmWWHa/m/74PQS4lzEoiROalc13NnGozup+y8HFnBjCNotynECViBKJqVcrMqaZlmVmKxzFhA4INRbhLXEKqodRptBErddxEEmftFZi4CYHT6uBGxOv6h/cYStUh9XAZti/wmEMVxDamgt94rgqAAyna9th3CEGp0uwe0FXKr8wbh+2i2VL+6BNpZCrSvBMtTQNn3Riun1Hz5jqBwiNEBfIfeUWM4nyVwbhid8VbDEuXiXfDRHcWGZeZeOC6m5eZ9YtS8y27/AMyMIv3g13BslwyzQlQOFys8BKeGMTkCBcquLgMui4Cm7qp8y50sTSAgZbVj2mLiAkvZEudM96Tfv6RK5X7xSuKGZYGkfMC4KmhXYu3bu4YqoD6EAKuCPiai+Wix/Q3HsiUY1Vku+6w75rFdUuY6w5Bq0R/gZnOs2e7f94GELNTfcrEvh1Lixa4GbORxLElxY7lUy37eibj9pfGZTAqGCdTqVccS88DLlVKsIxnG8wlVKrM+YRJ0EkEeVe/f9zMBPuvG+Xn7EqG0RQtMqVxWpcpH2Yln6UTX9BliknXBbJdioop1GajPgS2AK3+Lji35MVyXafVYe9RxMPBB+1f95bmCw+b/ANiDLh5l54J3wtMW5dMtgQJUqVKYlcLFj1xT9vRPhEjvhVkM8E0SpcWXTLIONzUHPBjc/iOIJO/QkG0yqlUC6Rb++8NHTjOp+FRRlebj9AfEUdMTwxct61ExuZK8CmxqrvcNR6mxGKfQWadIDMNAEIea6AX7TDzC37Of7m7gR5H+glLfZ7qrfYy/SbbwfUBS/SWDa+xUv8Q1wSotyoYiY4uHFQOD7yrnifMcTcup3OoD9vRw2LmECErE6nccy1iy4Yi3NJcGDjzBv3gkvgMWXF4MjUAalfX8iNP8kgCsGMvtB1Y0fSbNB2RX/mPdb6Rx5KiqOdxcS7MwqM7iAmM11LsMN3ZAS29+RKh2Ye66mXC5jY4IHSMGC+K/qMYF0T7f8gANn3AlWSoFRZRw6i4hublTUvgYtsHMZs4Tis5n7LwQzFojmDDioz8yokeM3DEu4NS/EuuFxSal0RMRai943hCEzdZHwb/iBRLHMFrH5mSGvKd4X+0jG9qC+SOH43NyX5EYuWOCoK7naCll5qEK7mfrT68f6Sv4rH6kfop+/wCsNfAQBTpHdr/uMqKhy8Ww1Oj9xP6hqHH0lZixfM3Nxly77gy79pqX783FjnhFn6rwQ1NpdzxwMuy+F+0X6xjMVFm5cGXF1LYMILS7mZfmFqrJjWx/H6RgyhZq5AIlCA8AQhXbognwwezLtrc4/wBiSyF0+sI4f5iiVdNXFpzHMOWGtxjLZQwvsKftKis4svJ7QXFPQFiaNblEc3GWL7vpMJjfavJ/ybJl4+SVY2QHgQf9wcweLixfvGY6jqdcVCa41Am59I7lUy88fsvBLuXTNS75GiXL94vvHLBuXmOpomowMGXBzLl1Bg43iM2unDED4Zf9+kDKGFdTftLzBIQhe0Z9Mx2HarEC1wBvYYz1EQE1juXblvrRyvqFIRKHx/0yoGqLSRre6Z4P7aHaLWmdeGyDqlMNW/Dh/mOO1I15njAv6WP9TTBqDLi8LCMZealVBKlZlcVRBeer4/VeCMSpdQcTCZRWXiN3C5iKxSMNQ8Qle/oqXBl4qWw1fvI/fiMKCtYaD9YucAH3Wn2HAvifCBATtIUGQEUuohfXhcBrL7jMBsWliWD3sr2YGO1IKGZbRoYtmr1LZS3G4ZoS1ZJbGQn0hFdoLGohisObmRlRx1lIB1e0IGlO1jecn1l+OxGUqz4i4nCn2my4e96pP4YZOGXUuL1L4trgMwLZpiF1xWJVcLjipTCfsvBL4uHF5l3mXxbMVH0BKjKxKqVUvPJLnsoOf36xAYAfP9gkA8SXXQB/DDKViENGBRLRaNsWD7ipVfo9q/mKrGwpE7GIiXxbvN41lbhvXtLo94VcTp+I1PaimVNs7fclCUG46sP7jVylN8JhDQRBQllaoJjFNF2VB4DXaI8jLdTH1mJ6qx7Yf3Bxccypd4rhmoYYN8GoMMxYuZeJfBYvF5leZ+y8EuXwTUuDmDLhNxuVDPxKJX2lSsQhMRLlQ4ILmgtlFzKHz+3KcVta9x4+hLaKUHulv5YQeGOTSV8ALM2FFJVU60bOpZf46yvD1Ktd5jPzllQzs5rDvxMe18GrGWvS2xta4t7pMMIWFGr22dQVSq4N5GBz9swY0PmtN/UUjsI8s9kVWcHYRdHbem5duQ5v2WyvipbxGy9v+uEIYwDKhpGCHkAj9OC3LnXNwcahLz4g1cuE741F1FnUWzh95+r8EWDB9oS8S5cWo8VCEMQc8XPwiw3KZvknkZKK955CtfG5nalyUWP8FCE0FB7SyoNQtw+SWSqwKdKZOyEQKrEI0ZUpUVfEV15Twzbld4DAbYwSBdQjFo6rtTfUIhaiX3cNOIqYaxKlNqvaSkC4veHmQEBGllPR7EcuJgQeAL0FRCOG7KqY3muvEcj5X2WG/hsgAAxC3aGLESVFGBaLTafWayLJrOiv6474L8TvUqI2zPUIp1Lonwl0y4t8DLuYuVepU/VeCXCaWHFy8RcSrlVOty53wc8XLi54uXXFTU/393X9xqIA6x+4i+0NH+0ZuOLly8QYVjaGhKwmigOwB4AfJcrKpANidRGWS+lq78y59x/JK2VH+kdxJWS4QXCCY8xTJf1ev9UxJaV8YH9wqyryYNJtfcSpnD13VWrv5IKkRYVizUEQ4sVgsfhINwzwko42MuoeZqajBl5l1UGLXLqXBufsvBNRQcQnvF+0I8L8y7gh7T6w9psmpfBhdQZdS4NEZTlgCBbsr7pEYHiXVM/ambooCMlK/sS45jNSrIrzLleKHlzdGWpSgt9slRSx4qt3iMBSKgZetiAUzxNMGh6NVgdXATOghf1JXygpGGW0bHhF8s2BzkhOVQJSKvAZZdMeYAUfZx/qKtVzHzTS+ajqJ9OIwH+oPyALPOpLLimTEW+hy+/5QcwalsuVwnAxYPDXLKuGJuVmG4YzP1XgiYvkwZeeL9ovBmD5huaKhEqamyLxc95pct4dRXlvrDPf4ISKG1BSjRpc+I4uyPulD+Gbj54rHANu1VkE00i/eEAgWGdC/oBFxzYuylyKpkbxTEfV2mhZSBgNaplIQhqzI56gydRX8YIG3S+CXWvtw1TV+8kLQhr9f9QDl+GZLgobWIojsuC9BQ7+a/uXdWNGXiKXMaVf9lROBL4HuO2DN8XBl3LzLt+IQv0JmXF1f+ZE4VNQzL8S+rlxthDUKjBg3Bi3Ny/aLcujhZudyLoeXqAGOFDQKmOy7+UgHlP1RLfys6hxdk+s2IaEUN138QY3dRabYDAtaDUzCRHCRIiWInB8fiAtcZqoMKj/ACIX6/sMCWqyEGRkhL0WNCkf+xK+gLKN5lzrvL71GYcwuCzN1ql/SOdsYfcz/UojjIxK5sFv6n/JeI4S7l/SZS+4vnhcYvgzAhKhCUqY58r/AMye4RHuLGGhLjBsnuH3h5D7z34wbJ7xAuyHmJ7hMmye4Q3WSzsj5SWZsj5yNTkmjJBuye8RMQmZfGf6hS022tsU2065xdPECoEnvEPIT3iYtkQ7I72JhaahfeEBKawyFZorNXRBqUoBBgB7NYN3mVN2F2TWKIM8Rq/+Ex/L5f8AUeyPl/qKMGqRSqw0gdwaIQbUPPvaj+EQy9fCOIU2zWEf1BDdK2xGcYMfMUzZ/hA1i18w1YD5en4iDZMmyddkPMfee4Rq2THsmLZPeJZ2T3rTBdkLNkOpJ7hB+yYN4RDVkEzce7GerJ75EDvX8RP/2Q==" }, {"x": 968,"y": 368,"w": 40,"h": 830, "type": "color", "background_color": "rgba(0,0,0,0.278169)", "border-radius": 0 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nMS9d5wlVZ02/lTd1D3Tk4cZGGSAgSGHIUdBQJegrnENGNbssoafq76GVd9l1113fdd1zeJiwiySFMkgSM6CxCEOyDAwuXumu2+sev+4/dR96ulTt3vQ9/MrPsO9fW/VOec53/R8v+dU3ejb3/72p/bYY48zy+VyrVqtIooitFottNttVCoVVCqV7H2z2USSJACAKIqQpikqlQqSJMnOS9MUALLzSqUSOp0OoihCqVQCgOxvHtVqFe12G0mSoN1uo1arodVqIUkScEztdhsAkKYpkiTJzuE44jjO+mi1WtkYW60WBgYGsr4ajQYAoFKpZOe2222USqUMS7lcnhZWxcnrkiRBmqYol8uFWDm+VqvVFysAtNttDAwMTMIKIBtnFEUZ1lqtlvVXhDWOY1Sr1aytdruNTqeTw1oul7NXYtpWrLVaDc1m8y+KlX871mazmY2lXC6j3W5n7bAv9hfCSl0lpk6nk80N5a7zkiRJdn0URTmsvKbT6aDT6aBSqSCOY3Q6ncw+Wq0WBgcHC7Hq5+12G9VqNdNx6iaxdjqdTA94HsfYbrezOUrTFKVSCVEUZX2x/X5YW61W45FHHvl8dN111zX233//apIkk4w6iqJJk9LpdDJF4SB4HQfACYvjOBs4D7ajwlKjK5VKufPZLgXMzzqdTiZcfs+JA5D7TJWS10wHq06e9kvFIw7HyjaKsPI79s2/qQzsrx9W/k2s/I5CV6wUPhWlH1YdNw2G43CsKlPFrfPA/mmQnIOicRRh1TlyrNSR6WJttVqZs0ySBKVSKcPFw9v+S2DltS5Xxz4VVm1LdfwvgVX1WvX+wQcfbMRRFFW1AzVudQgAMuXxCFIul3NGp0bBQag3ppHSsDkhnDAdaKfTQaPRyM5RgGzTjZDnlUqlzAvrBOhk9sNKpVUBEatOqkYAVRp+p4at7THS8DNGCB9LCKt+pwJX2fC9zonOdwirzku5XM7kolgZsdgWxxTHcRZItH+NqvqdsjfHqoZF2SrWTqeTi5rTwUqnyIipBulYVS/ImImV12k7/bAmSYJWq5ULeC5XnQd3RsRKHP3s1bGq86GMi+RKJuTMaQJrrVypVCZNshsdB8+BaTqhXpWTF0VRLsprBNTIyXYUMIWnAqNxKiNwQ+X3nBwaQLVazQlIsYYYAA9OrGPlRBIrz1WsIZagiu6KGsKqyuZYPeLyfaVSyeTF893xeH+OlUpWhJUUX41HHb1G4m3F6obeD6tGb2+/CCsdYIiFdTqd3Bw4Vu1HA6ZGdB2zByPHpayNx1RYtX3FWsTQ1HGTUQDIMOn8U89DgS6TK3NI7YiDUeXXi9XAmI+xUVUyTmTI07s3Vk8X+syF5RRPHQgnR4Xs3pfjV/bAiWI7LxSrshjHGsLGv9U5q5NxrKp8LhPFqornSq7jVqz8jFjdYDTNc8rKMSnWUqk0bayagm4rVkZRnh/C6rpBrBwjA5zKtR9WZcKKS8etf6s9TQerOlteS2euOuyOWBmXprrEqnUdbVv1xLFOXFfOOvZoyUGrw2Ckceqkisf2lGbRwHQCSPF0sgjKGYOzCT1Xr9G/VSAqYI2WGs3UKWkk7YdVjWBbsXqKo1h1TBqhvF89350Ax+5y9Ug4lVx9LEVY2Z5jVYf752INYQCQ1ZZU5ho5i7CqU3CsbLcIK69X5+hYdR5pGy9ErhrQHKuyO2c0LLCGsNLG2S8ZjGLluDqdDspuHGqIPDx31yKXRyZ6W/W6ToX0GmcGCpIeU8eizoveUQXqhu9pi2JVvPo3cQCYVORSJ6RCdMwvBCuv1f5pvMSqhuqK7UWq0Ny5Q9foVISVh45Tx+tFMzon/q3zxfNUN5QCM+rq3ClWvur3RVj9vRpWqKDXDytrHY5VmZu3wfPcMStWTyn6yZX4twWrpsj6vY7T6xOKVVdw4pBH8snv5ylpkKrgUdRbflXl0+juVCdN09w1mmN52wCyCrAWD3VZSOlYCKPSOPbv3p2HCoa5rbbHZToVgmJ1NsGxKVYKVB2GGl8RVo4jhNUZHvv3/Fqdns43seq5xEpFVKwqH438Pj/qWHWsEwqZc8g6pyGsilHTPo5Z2UcRVs67z32n08mw6pKpswPHyiVUl6ti1fFrmq5YdY54nqfRIQfkWFWP2aYvLrDgrFg9dS5rzsVJbLVauZxPwegAne5r47VaLQdCaap7SU4mJ4oemW1pgYfXsV2dVFWcKIpyS4HeL8faD6viVawqfAC5ImoRVhVcCKsKWPv0/JrOSZUKQBCrKn0RVg8E6kCng1XH2w8rHY0aGp1gP6xeCCySq1PnflhdVkVYWTDWeQlhpT0wIk8HqzLEIqxAvuag41Xb2Rasqns8n8zVC+TulGKfCFVAAtcJY7T3hpwtaKFIgamh0wPrhKvz0ciggtIJ0InwiMioEGIJ08FKDB6tiEOFPF2s2lY/rJomOFaNukVY9VpXbF06K8Kqc61YGb18XhQrx+JO07Gq3hRhDbGiEFYNBDrPjpVtqHNyh+UsMDQf/J7L1c5evV7mWBWjYtW/kyTJsXZ3VMpQ/lysoaCqWCf6mZwisBHPoeM4znk6HUDIELTa6rQvjuOs4q5Gzp1rXApM0256wlUbLSqp8ulY3RBd4ZV9hLDyfMeqOLw4NF2s6uEdK5WPdNCxarR2Z+DFLk9HeI7mvEVYi6IbD+62LcLKfNexsi3KVanvtmLVsbpToq4WYfW5UTk6dmJ19qXzRtkRq26K0/SF+0oUm7NrbV/Hw/YVq56jTqifHihWJwiaYvPQIFn2AYWEooNVgXAQjHbqLLjO617ZDzVEnsPJ1kGrF2RRUw/1slo8YjTUCVNl1EigY1Ivq5NKrPrZn4tVx8oIQUyK1Y1fx+Q5ahFWtus4VZlC7fIfqbbO6VRYnW2q0jpW/j0VVr53w3WsvtTqhuMyVGfjexVUH7cFKw1R26dTVMbWD6s6glKpVIhVZVIkV45F0xJN41VHeEykKr0lRG1QjZ5CZcda5+Dg6TE1X9N2G40Goqi3fq8ToAJygyMQLRb12zqsCudC1qowD+2LwiBWLbJOFyuZUJqmOazs35mJUz7OMdtSrEpDOYZtxarz7ljdmIuw6ryRhvP+E35ehFWNVfsiFsWoWNkHz1WjCgWXflQ8tELAPRZTYeX26W3FqlFeAw4xUv4cg8rVA7MzAh6OlW1qGsTAqFh9xZDtNJvN7F6TUqmEWCl8SFikWVRAKpgqFKkXB8Abd5ReDQwM5NIOKq22xS2xqtQ0OvXEBE9QOmZSXPewnDg1QsfKdIFjptBCWNk3d8Bqrskb8EJMiwqjKz+O1ZkCsWpFPYqibM//tmDlOSGsZIeqZMRKY6UhcUzlcjl38xL1qQiry16VXym0Y63Vajmszip0jouwqjH6UvZ0sJZKJdRqtRxW1RFi1bFTJ5R5Ola9TcDlyuvpGByrHmoDxEobdtZCXL4krAF4YGAg78x1/zhzaFU6DozelwAZdZRlKBCNWjzHvWDIcbgX1CKPMhtVagImvdPvPHKzrxeCVdMbp8Kam4awesHL6a1GqX5Y1SBCKyn9sHok4/VFWD1Pphx9NcKZYhHW0LkhrPxb+58O1jiOtwmrM0KN/iEWq+MP6fB0sYb0tAirOogQVp6jjtSzgSKsmm4pVo7ZmVpMkBQyvZtGGZ7MQwshoc1GpDDsUPNQvY6enA6rKB8tlUoZ9WOUYBs6KcRAg+NYdYLofLYFq691q4dO0zSH1fNQp32a81OAqkiOVfdYKFZNzYqwauSgY1LjVxycc8WqVJbnNxqNnGGpQajyhbCGxtgPqy7x9cOqacILxarGwzb7YWX7tJ0QVneGTNVY+GR/ijmEVdklsbZarZwjUwwqM35PrOyf54SwqoPSQFpW76SRLlRc0bxMz1fvynMGBgZyBRil1uoE1AB0l6IC5+SoV+Uk8hwtMqpieirg3pTteMRwrG6EqiyKVaOKYmX7+syM6WDlHL0QrLze0x3PT1XBXK5kCcQ6ODiYYx7anjqM6WAlbZ8OVp1Dx8rj/w+sbI/PZGHtQzHyVetbLxQrXzmnqpvan7NWYmLbqj/ESjvlebw+030twqnnVaWjN9KI6SB1QnRieI2uNqhh8mg2mzn6pYpAdsJoQE9O5VNhaiqguNSAVVnYF70vlUaVQp2eYwXy26zVc/ucsg0Wyrx/nq8pHmskxOpMRNNAvmodIDTf6rxDWJ3OKi0PYVVWuS1Ygd5qRRFWRlhPeTkuT/t8mVfTqRBW7WcqrKrPjpX9cD+NYmV/xEosaiMAJmFVu9HAo1h1LlV+KpvpYg2xY/0Xa5TXnItKR0+nDISTo5GEQvNlvlDK4hFB+wl5ZG1DJ4yFM3VoHINHd09rNLfmJIaw6rXqnBwrha1CdoUi1hC95z8qjEevZrOZKZhiZeFPI6VGIUY6NyL+7RucdEWEWHVu9Dzdru6Hs1OVp2PVa4hV01PFynlzPXJmqm3ybzUIYtBawZ+DVWWlWENptWLl/DebzZyBa0HX2YNj9f4YyDygK1a2p8u5lFkR1tipB6OrCkQnUL2SRnKNEPxcKSZB8nql7ZwkvZ7fRVGU24aqBaRKpZJV47WyTrBqeBqVef10sKrwXyhWxUMKyPYdq+ahipW5PbFybIzayvZUGTgGj1Q6hxphPPXUXJpj1SJiEVbOrS53hrAq61OsUdRdFeBKGJ0Ir1f25FipW16c1CJ4CKvXVRSrn+tYqacui9BKozsmOodqtTptrGo/QH5beD+soaxAsXJ8jhVAd1OWd6QnqQfXiEdaxclRw+JnXqjSieKhexkIiucpLVOPqMA5Rvan/erkeL0jNPFOlT16ceyOVaOVzokWUfkdPbxj1dRCsSp1nQorDcaZi7bvKZpi9Zy+CGto2VGxauSbDlbd6+HKrG37nhPFmlFl0a/QjYw6hyGsmmooVj1PUz3HynFSb9Rxh7CqbennXrz0+4HobDXI98Oq+uRY1RZdZ1ResRf7XPlVCVVBtGLrCsHvFbD3QaPRSVWFo5fjdb7dm0BI/b1wlKa9+1g4VqfpTh+LsKoChrA6I/C7ZZkqqeNRrLq+T6ycH3V2pIiOlYZBxVWsmi72w0oHVYTVlVT7VaXWcU+FlXPlWKkfilVZG6/1YqIySR0vx6d4vHCtDFT1VLEyPVWs6vyByZsXlX0qVo5Hg61i9fRBsTprVqzK3hQrD45F5TodrHEcI+YAlMKpN9HGtDP1bBwQAROgFrbUuJIkyZaRqEwqLE0PdMA6MVpn0POUDmtBh+8pAMeq1xVh1QIo33OeOLnEqorAdElZnGJVwalwHKuma067Q1jZv+Kiw/HoqpEohFUdbRFWVvOLsLrz0e/4XnVCsaoDK5KrpwcAJmFVQ/MApVjZr9Z09Fxi9WV87UP1PuSMlAEqGwnJ1XcKO1aeoxhCWHm+b9mfCmuOWbggSUlokBqZ1Eh8lUOpsdM1fqYPq1GmormmUndOptNOjZwa0T1/Dq3kOFZO5HSwKp1W2uYR3HN2NQjF6nM+FVYawVRYVa46z1QUff6qzs//K6xKcznOEFbqhjIzYlVdKpKrskLWPFgH0cDjWDV48Bw1bseqzrgfVjr/EFb2S1vgI/19WZT96fwoVo6p3W5Pwkobd51W++TnGih1DoGJAieLZjopSg15X0eIyiq99IjHQyMY21dlU2+pToSToamGK4MvU9JphJwZgGwrto5Fz6/X6zl8qjDKFoqwqqfnqzpMxRjCSpajbEsd53Sx0vHp8yeUCgPA+Ph4X6xUJh2ry3A6WD1d1TZCWEPOSseu3+v5+gwVtk2jGxsbC2LlearPHKtG7xDWUArkKRz7AnrPCXXnrFh9KZkpiDLDOI5zWNk/2YdjVd3RcWmK5ONWdsZzYn0+H0/WTrhvnKAVrE4i6U+ocKKTr55Xz6HS+CRSWYA8pVOqxevoUZUK61g9OqtX5ZhUMEpxFavXStzY3ZEoVjo/xaoGoefxO3WUvI77YzTFCclFlUCxxnGcuwdBsarMKAPdc8DrHSuV3bHq8hyv5fc8VEYh9hHCSlzTxcrPFatGUnVK6jg9LWdg1LoHdcJZg6dcRViJi/bG11CapRiVYfCo1WpBrCpb9uurPZoaq1zjOEbcaDRyXlEnUdMKUqRQbk8j1BtqeCid05zJo5RPiue4HhFUyPzna8vq0XmdL69p+8RaKpWCWHkOz3OsSudC+bZi9VqCOqLQ/On1bNOLxsTK6/jesSoNVaw6DndU7txDWNmXG2Aov1ZsIcNiW45V9U7rAp6WhbCWy+VpYdU02LHqGB2rpiFuoO4gHatGea0JOXNRrL6KqAEnhFXlwXH6XiHHmnNsXlBSwH6noHt1Ba1Ood1u5wBp9NH+eI0bHo1SQapDYP9eHKTi6kS7MvNz9qlUWfsLYVVBc7zEyveKVff/O1aOOeRM+mHVOfJ6kX+mzGs6WEPUWR1FP6w8Rx1ACKse6mD6yZW6pzINYeV5jlXnVbE6u1D9CWHVFFFlqnPkTkAdJPvV+oE6AZ6nBqxzqePkeYrV9cixukPgnCZJbzHCsar9ZHedcuAUFgtgSrV1QF4I4oBckM4EnM6qIDWCK01T5VHD10jPa5RB0HHxmmazmbt9lxPlWDXdUW8cwgpMXs0JMRrPf/V8bU+XBf3OVDd0xco0kM6e9yn0w0o5OVYfm6dBIayuF/qZt8fzFKt+5/PHthyr3gJA3fCag1b9Q1h93LrCojqh54SwulNQ5+tYdW54rm7qC2ElNmLRDXuOVesc2l4RVtf/IqwxG6VHUWMPUe/QyoErhuc6BKROQj2750geibxuok6ISqPKQnCqoFHUe06AYqUBKFY6mJxXDWDV6KXtOVZ+71h1u65i1WKzYtVb8R2rCjiOeysTTM10hUodst6LQayai6vC9cPKI1RDIG7tl1j9iWccowaxEFYakaYNuvU/U3CZ3yKsGhx03GTHHLcWNHmeO0aVsbM33YmsLEGZmQbDEFaOV7Fq6qCOVm3ZsXIc08UKoHuLOidQBwd0ix90Dmp06ul4cGnH6bZPmgKjYvkEUeF5DYWik8z33CLL83xVR52XY2XfipWOKYSVfevautJQ71cppGJVo/B0y2lqCCuVM4RV83s1DD2fUYxYQxFIaX0Iq46tSK7uUEJY/X4N1Scdl2OlThRhpWFOhVWNIoRVDVBlwe+VpTjGIqxqsJoOcFwhXVIdVjm4XNmet6FY1XFMF2uSJIjdCDnxTosVjP6yuCqFOx2dEG+LNE/71HNCrERTE1VEZR1UIGcgZFCKVZWbfasDdKy+fOuRy7Fq1FGsodREaZ/ing5WbZcOT4XN7zhOpaHalq4ETYXV06AQVneWGk2VrTpWjufPwerzWoSV41esHqXdGYQcNs8NYSU+xco+piNXtluUwqiM1Klo23QQoW3j08E6cV6vAy1uuIPwyQ45BvWYQK/2kct7RDi+CqNAeD77VA+rdJiKrZFb+1ChaFrA3WqeczqLUaw6Ni+ahrAqfSzCqoxKDboIq47PGZ8qTBFWj3rqoPhKQ9wWrBq5+mFVZXSsbLufXEORXbGqDnukD2ENyVUPjsFvVw+xJKBH/6fCqvPUD6satUd6vQWCuhvCqrYQKhSrnRdhBdBdDeGE6f5zFwwb1UlRFqAdagTjgNRoqDiag5FpaGTVft1peHTiJDBH17yO12pRT4t8HlX4vgirOpZtwarpj/5epfetWFW52Y5iDUVPNdw4jnNYQwzSsbIvxwqgEKti0dUCl6tjVcelbRVh5Vh1iVix+v0iypJDWENyVX1Wyq/jC7HpJEmyuti2YlVDVqx0tkVYndGqPmggcaxsR5k0+6CDmBSIOLBOpxMUFkFqBORA1WvSM3IAClaBeqHSaR2NPE17z470/t3LqlBc4BqN+bljZbuuKIpVnaZHeo1uSm0dq1JEYmV0mA5WF6oaso+H/XF+FauOR9uLomhSCqFy1aioGBxrSCEp1xeKVaOnGkQRVm1H9QLIb2zj9xp8tL2iABDCCvRSVceq860R3V8dq8raxxYqQjpzdKyh9lSWxKByYx9l/dAPBaLUSj0dFUnvC9BOtV09XxXXjU330GuBkUKh9w4pUKiAyOt0GU2dgzucEFalnlp8c6whr/5CsALI9vmHFEWxKjXdFqxUJs4h+yjCqk5CKWo/rPp+Kqz6IGCVq45jOljVuN1wtF2Oidd6pOa5nBN3uo5PxzZdrNpPCCv7IdbQ0nWRg1R5cEyUs2J1mXPMk5wcJzu0+5GKyQHx0E74N2mOX6fCD1VzFZhGM062CoQT6Y8u46S5QSmd4+TohCkzUSMIYVUF1rlyrJwDXYriipI6o5BiuQMKYQ0xqKmwhlIQxeoYFStZmPbF99uKVQ2beqFYPQprVOP5jpU6RMyqY0VYPfpSDlNhJWOgjEJY2bcap+JxrM5gHKs6EV25AMK35HsA5Wf+SqzaVwgrx52mKcr6UFUFpfmvKpFerBPAwfMI0Rh1HkqRCI5tcKD0dk439YlCakRquMoQ9BzNrZ3O/rlYVXk1Smqf6ow0n9xWrOoAQljZfj+sPF4IVqBX+FSsdAjqIG699dZs3Ntvvz2WLVuW9atKqvdv6Jj9yWehlEGdQ7PZzBk258BrVEwTlI1qcVYZTLlczgychdQei06Rpr16D+ed4+A1ii2OYzQajey9snBlCWozztZ0Pwn7VRapbCt0nQZ3tR/6BMqDc1VWT8rG+M+XepS+aETh56ogSlMdJP+Nj49nP1DjVFDpPMfoy2zOhHSi1Mur0qkRaLRVo+JEKh0swurUXQ9VjBBWLX6GsLI/x6rfOxZ39kVY1WltK1ZXPh1bqVRCvV7Pis5JkmR3QbKvUEByZqgOgzqxdevWHItxJ9HvcDasOjnV56G/VU9azQbK5QpK5fyPa7O9osO/q1QqmD17dk4nVK7qvNyhUJ/0OrcDlasGan6mxU13IqVSqbsa4jQnRGWAfGGEDfBzVTw1XC9E8Wi32xgYGMgZv95LoVFSn/mgwtT80VdmNKfl39l9+XF+PV+9N/tQx9QPKz/T8SjeKOpu5Z0Kq7Itj/qOVY1K58nzUyqL1lI0grxQrDpudZBx3C3Y1mq1HLNUqu79cGzEwLZdBxWrHqHvQufxUCf0Qg91fJ12G1EcoVQOP4y636Fj93+e0gN5I+c8eQ1F56KfvXpqpu2yL3VG7XYbZVXsUDRSZeB5pGQsvind9kG6QbgihIqJ7Jv/eE8Hr+EksuBDhVc6z7+dljn1dUeo3lTpp1aTlQI7Vk8XlJX1w0oj9D0JipXnhJbxQlg51v+XWJXZaRVd5yEUdHi+6oOer9HSC+U6b0WHGq2OcapjOk4nc7BJgrQUo1yu5WTm7U2X/QCTmaTrw3R1WN/TFlSuXg/0sav80nTiprUQII0C2pgqI/Ma5m8axTSC8u/Q7dIKjOc5PfJ+1blRkTRfC02e9+fKo5OlLIGfk6J3Or0NThoRtTbjdC/U/nSw8nrFSpxOE/l9P6zOzBwrr9FCYQirOi1idaaikY1Y3dhdDhqoaCy+bOsOytsrYh+OW8/nd95myOj9KJXLqFZrk6Ky6+m2sA21NeqIp6DaXj+5apt+h6ler46bnzlTj6Kot91bI5NGEy9mAch+r0M7VE+ngw/dyMT2NIUgNddqthZstNDk0VAnRR1dyFg4fnUGjlW98lRYnenoOrxT9uliZbshrCGnzrH3w6rthrDy3JDR6rWasvDGNiqoBxliVd1xrDyPqaZGQ68vqX7xKIrm7hiKvi9yMB5Z3RkUOa8sDe2En2sxnUPbDcmVTtpTO/bvGPQB0Pw8JFfKnkVfDWjtdhtlCpMdqcCA/I+rcolVo48K1FMM0jWNDF6B5fX8vVCl4/RwIe/Jw5cFNaoRsBZcdZwa+V4oVo6xH1a9pgirr23r3hLiKsLK80NYdS9EiEFo9FL2osqmyqo1KWINFXcVqyo251Gx6nIqxxcyUD+2xRDdcUw3NShioaH2NaonUfEGuH59q/6oc/ZFA90BHJIrkHcuzlJ1W7rKJU17TFp1MI7jLrPQgTYajUnRiJREn0akwmeHunasqwu64qLRkkrDaryyCE+DdCJV8FRaPWh4pMhFD3dpNpvZ8pZjJVXrh5Vj1WXnbcGqkcONLRQVi7AyyivT0us5Xj5LlYfKla9OpVkPKcKq+DTl4PwrG1IjCNFqx+qHfh9iCzymm6YUOSNvO+Qw+vVN5qhsKzSWfgfx95MrAxafpcrPNVsIyZWOgnJVx6BBTmuOE2PqrWMnSZIt71EZQkxAUwxNK3S1ged7hGAerHmeDkwVT41Uo50bjQuDqYAvhzpW/hwBJ5h4tAahNRfHyu9DeXUIa8hBKFa25dRzulh1/lzofE4GFZUBoQgrccRxnJNrqF7CcWjBmbiKag5Kn7WvEBPzo8hRFDkCnbd+Ud0DUb9+p9POdNmLH8qsXa7A5GeN8pmbAHKOnfNJHdeHMalctX3VPepQttwdRVFu44/+HF4URZOMgo3EcYyBgYGcUnAytfqtikHw7tU8T1aHAfT2BbD+4aDVm3qEU3aSpvlNTuocgN7zCD0loEB0HZsKoXNShFWLRf2wqmPZVqzOTkgnFas6EH0mx3SwqpIqXg0ijlUjWoiB8Dru/tXdkWoYaij9GMJUxqlj4XhC7fVr06/ZFufSz+l7e7qJz1mnblH3Yro+CMoDfa1WCz5WMMToeI0ub2e/dUoB6qYrFkZUsARCxWfVWiOF1wJCVX0tjPlGG6BXlFHHxTH4bkc3VB5Kg9Ubq2Gybf4Yr9ZaVGghpqVRvB/W0O7NflgpNArKHYRfD/SKhKoImvNqvabRaOTkVoRVWYFiVTaoShVScjcYvS2AfSlWYvEIp5FalbwfpS9yAtM5QuxlOowm9Lf2604j5Pj0O5Ur0CugegGSOsxrVCbK0Mh2fZzuQFUPM3YaGjw7qWP3CMgAACAASURBVNVqOWXVDngdqadGaN3o4dFEK+GMRLVaLUdhgR6boAPz/hWIfuYUXh+Rp2N0rAMDA5MYlGJl2yGs7EsNRyebr0x9irDyvQpMI7IbjTtRxxpqI4RV2+yHVc8NYVW5MCD4d5oeKnvQcaqTdCNxRXcHws+KHEi/w6/z996X200/RzSVQ3EdBnq3+rdaraxmoYsRLgfOpxaMQ2NUm3LHS32iXDW4xdoADy3SsZCnTsWjtFbQnZbTK2qbmgepZ2RF1tvUZyw4u3HnRRqmkZoYPVI6Vr1BaSqs6kDZv/etEdojqGPlfDhjCmFVpWBbLnB3isTA9743ZjpYtX/tWx2Tjl1lrxFKsSpzVWMIYVU8Rf/02qkMVFmSO8t+14cclLcbOkLnhxwPH4unjFuDID9TnNQBzqnKNWTjLld10gw8KtdSqdS7RV2ZgAuYdQyN2LqfgG1QiXi9G1Sj0ch+SUlZhralA3dvHsrDPNqxTV6vaZVTao5dsWpxL4RVDSRE+6eLVR2AYqVAi7Cq8Fmk9EJWEVZN+fw9X52tTAdrvV7PYeUYyHQ0GlIhXwhWVXKAOCf/HMB0/vZ58vNChu2fu/Fqu36oYWu/oTZcrn6+swDKkjrGVE+XUfvJVeWmOqNyTZKJZ3CWSr2nZAH55ULSSfdUHIhGnNAkKNiBgYEcY4iiKFu6pBejk+FYtEimqyIaeVQBvRCmHpnvlR4rVuLqh9XZhCsP/w0ODubOj+M4dxci+1asvkyrWJUFkI2pg3Uq71jJnDgWNVzFqoY9FVZe51hVroqH8iRWnktF50Gld6xJJ0G71UTS6SBNUkRR3phChzsIZSD8rN+1aZoC2fnF+ytC/ek52/JZ0bYDHa+fo8GUDlprFcrsXK6OmUFH5ZrVLFTIbJiT4LsIeQ5pitJoHh4p+Urqq9/zJwfZnvanqxXq1NzQPZ9nH36XKZD3sMTKSdc6yXSwaqHJ+9dlU8XKcatX1z6KsPJzxapGr1idZSlOZZHOzEJYda6Vpamya1QLYVUnpEVlHQtloI5PHWvPmVcRxZOXYP3QSB/6PPRd7+8Uq1c/i5UPP4yN69eh1WpO9FnCrFmzsXzPPbFs111Rsh21frhTUhz9DpWvBhA6Xeq8zh378GK6BiaVK52Msma2wfGpXLM0hIdu8NEbt6goGplUkbVARxDsWBmKKrFHRTVgjYrqzHg++9Anb3s/ACZRZ1UgGjGLR+qg/lJYicWNQbHy76mw6hi0H83pQ1jJDPth1bqBPsOS86DKqU5RsaqTLsKqehaKcurYVGmp+KVyCYh68+IOWo+pDNIP6uGDDzyAm268Hgvnz8WSJYuxx25LkSZtRHEJcamE0dFR3H37zbj6ysuxz7774+hjjsk5fY63qH/FVPS5zonLVZ2+P/BH2bkGPrbjcnWZKlt3xt1ut7u/SMbOqdhuhKo0ruQKDMg/r4Cda1TSlMOjuyuJRhidVFJcOjcFx/dU3JCTInjFqh5UU58irFRg7QfoPQpPnYsaVIi9+bzp0Wg0gljZdhFWlQEVQ7GSqqpcPaJ5akAF5fW881hTLXUQygrYBrHqwWuazWZGg6nwOo9e6NXDDbRfesHv9X29Xsevzv0FKlGKow9fgScffxS33nAdhke2YrzeQJoAlUoJ8+bMwtJddsb++yzHxg3P43v/8x285vV/g0WLFvUdT2h8oc+JW/VBmZjan27cUpbgK1RFcuVc+t3azWYzt9GLjrmsikWB0ujc89PotSOnuuqdeK0/Acn3KlAJHIjmrDppusuU/fmSklIrp7J/CayqiGoY+gvWQP7R8OqsQli17qJYnVL3w6o4dbwuFzXYEFZVZnVwyjIcq6+MECujosqe7REH0PvxpiKs28IeoiiaKDGkSFGcljD4fOdb38QhB+2Hsa0juOD88/DU6nUYq7cmrka3rQjAM2vxx5WrsMN2f8SKAw/APnsuw09+9AP87TvfgwULFkzSC3cYOoaQM1On72klv+PcagDzpU7Oe2ibOA/XZZWrOqqMufjefY1ObIgD54D0O1Vyj3gaSdi2vlfnwsFyErh8pOPyqOKbe5yVcAxOdfUcx6qFtSKsRdFdsdIh8DWkOFq864eVc7utWGmsjlVlyv7dGLVIpjT3hWKlYrJddWiO1SOofh9yYiGDBLpuIqtCFDCSNE3xs5/8GHst3xXPr1mNSy+/Cg89/izG601AHQXbB9Bsd7BqzXpcfs31uP+++3DIgfvhB987O7fhyQ9lW8riHFdIrrr8nqbppFoWrwvJ1fugTP2uZ51nlSvrjAC6qyEuII+4KgRXLC1CeT6vCqGfaaVWqbBOCsehntMfudfP0WnNgcBDyuVY9bwirJx0j5CKlYLzzTJ6b4r2p1gpzKmwaprh41OD1T44Ls+BFasrtO6FCVXVNZhklFWw6rxwzpXROladW56v8nGjcpkqZh7qXPSclStXYmTTBlQrJdx40y1Yu2EYEVIkaX7tg++TicWRGECr3cGd99yHNc+uxsL5c3HLLbfkxlbknDxN0++UnWkqonLV+dDPXYfVSavs2b4yRdcLHpRpkiTdh9+oo9CB0Yup4in1LcpRPRoDk5c9Q8qr3ykYXg/0DI7Kyu99DBq9dDKcyUyFVdlESAjTwcq2eJ6nH9oPz+V4+mFVgTprcMffajZQb7RybQNAY3wM9WarECvSFM1WO4cFAJJOG2Pj9UlRT2WlrITjdnnoeJQduaHra5EhujxCn/vfv7/uOqw4cH/cfsedWLdxBNHEw3eBqPuadtlE9/MJRwUgAZCkKRqNFu6+517stuuuuP22W3NROSQrH5dj05pVzlBlzjivnrbSsWvbWsvzvUueBgK9zW+OI47j7o1kIe/PQxWbg1d6C/TWznUASlfdM2q7Xuzi99znrktBrVYLzWYztz9AnYtGqxwdFc/ruPph9bVqYlXv7hPbD6v3yfGTvqritNvtbcKqn+ewJi2c9/2v4LijDsNBhx2LP6zaBABo1bfih1/7Vxx52ME48rhT8OTGZg7r1s3rcfG55+Dtb3wVjj3pNdjcmajBNOu47Jdn46UvPgoHHXoUfnfPqpyTUqzObDh/Iazc+BfCGpIV2w05Af3nepCn5cD6tc8hSTr40+o1XVlmjCJFKQLiCIgioFqKMadWRinqOo90gmGkSLFh4zA2btqA+vgYRkdHC/v0f/xeD2fhrkPKCkIpvQcnfeCyO3O1r5AOazAH0C1w8gN6ITVQHko9K5XKpD0MXoNQQfl7tudKzsGnaW9Z1D0p23BwvJZj5DX0lLp/oAirK32n08n9crl+HmJD7iTUcEMKREagWNmG5pshrFpIVKx0qnEco9PYgn/+6Pvx3d/cgmMO2w+P33gX1m0aQ2NhBx8/45248ObHcNCeS3DbPU9iw+Yx7L5dDX+8/Uace+4vcfElV2LN5joWzZ2BEWyPOE2AThNf+swH8LWfX4VjjzwID1x3K9asG8kpokdSjjG0z8KxhpTWv5/OoePpd1271US73cLmTZswNjqGTspiKDBUibG1mSCJIkQAZg1WMGvmAEaeH0EcddMRoOtcmq02RjYPo1zuLq3Onj17EoPQo2hM1EfFr4xPgwoxUu5qf2qXfKYqz/U9OW7HqsPu1GJSP6WIPClEpVnQc7rkm5N4neetSonUM3KguuEJ6CoP7whVAThl1zGrkulTqThhPiFsxyMjx6hC1sKrT3AoR6cCcJyOVT/rdDqTHm1XhJV/K1ZeG8cx0s4YPvSW1+Fn1z6Kb333uxh55jEc/NLXInn6Rrz61JNx1f3D+MH3voV1Tz2J4191Op657Xy85IhD8LJXvhFX3/EY3vbBT+MP996DF++zPfY/8nA8eP0leOMrT8G3zr8VX/rW2cDmZ7H8sJOwsL0K5/3iJ9l86o5RjYauS8SqrLQfVmcRRe/1CF+TZq+YYDVduXWZQpR22cSyHWYjjrsfpmmKGTNqKFcrQBShM3FOt9Gu42h1Omi3Wiibbkz3mGSYxiC4vMm50/OA/C0XbEdX4qgjdC7OSHm9PjrCGXSZS3M6QB46EP6tUUIb1ghApdE9HGw/jnu/dMTzdV1Yval6UR5ecFWwNBQt8nAnIQ/FqmNXrB7VGK0dKw96a8XK6/SGLeILRQ7Ou6YxIazKJBwrN9KlaQpEMfY45Fi861/fieF7z8PdT67HwJpf4723XIGDDj0Cv/rP/8IDv/0KHlu7Bc/89hzccfUsHHP8CfjCdz6Mg/fZHZVSjJFnH8Lv73gYo6Wn8erLfor9Dz0aP/3VWRhYexOuu+dJVAbW4D1/dzM+/JGP5DZ3hbCGHLTLwOsyjtXlmGG1Q9mdn5N2fQSAiRu2KlVESFEpl4BGG+nEObPnzMbg86PYUu/KfWCghgQTTCiKMK8WY0N9YkUsjlEulVFvtDBr9mxwnbU3jnSi3/BmLR2vPsqR+EMbrDTAU+98jtUeyUyok9Rb1WH2qbaoz0Qp84d5VcActEYEL6YoQ6DCajHF26RCcDJI57USzsMLYDx8+VBTGR17iIZqROMksR99apS20w+rb4v2a5T26Xt3fqGag0YZHYNe6+nTJKzxAD78yc+iVCphTeVEvPlNT2DF0Sfh5JNejB0XLQSQYuDYU/Gm0+s4+iUn4+STjsP82TNyivb4PbdifT3Ccaeeho/9w4dw2P7LEUcRNq5O8dbT34zlBx2Nl5/yMuy4eP6kyOcrKByX1iRU0aeLVXH6ex6eAhSlBFEE7LHnXtg6uhlDM2dieLQBsCYRlzB7aCBzFrVqBaON7vt5M8qYP6OMDfVxAMDQzEG0O20s3XmX3A110hPyayuTx8vzFas7SOo8d+J6iuLPi9V51rlnW7qjlzLQlSjV21KphOimm25K99xzz0leX0GoMZCK09iVNrqQ+eoRgoNXUD4hng55u1pH4KFj1DaA/CPs3SsrRdM21Tu/UKz8TPsP1TSmg1X7UawUsmJ1x660crpYm2PDWPnUWuy75+6I48m7T4uw+vz87ne/y/paunQpdt9999w4nU2oo9RAMjw8nDG1otRD9SHkJFy/n3/+eZz1za9i8fw5uOn2e9DqdDBUjbHX8p2wdXQcDz25DilSHLL3i7BhZByrVm/AIbvOw5pNdazZPI5yKcJ+e+2O8VaCd73n/Vi6dOkEcylejeF7H1+lUsHcuXNz56jOcn59ty51RPdOsP2/hL0CwCOPPNJ9noX+88gH5BUxRK2ZlyswpTSsi3AAoWsYuXUjkBu0RyLdehyaQI5BaZ7mwuxXUw9PCZxa98NKQ1OsSh3ZfgirKkgRVhq0Y1XjZd86NmdhvEbZTAhrbeZcHLDPHiiV8u1xvHqjkWLVFRzOcUjp3TloCscxO9aQoRUxB3cqoUC4aNEiHHv8idg0shXLlu6ACBEWzJ6BcgTMmzMTZASVMscB7LBwCJvHWkAE7LjDInQQ4dDDj8TSpTshxCDcsakc/HNPxTjPKiev5zi71gBA2ahecF51Fyj1p59cYzcWjUCqvCGAHJRWsJUqseCnuxPV6BQUqT2vKZfLWfVXJ5DXs00tqOl3bM+Vg9g07dDJV4/rRdUirFz603HpeJw5hbBSITQy+PWKVVcXFKuzln5Y1WE6VkYrdzjEyojFNnWsni5wFyLHq87GlZyv/lMFblhTGaAa02TDAtSoTzzxJOy1/0FAHGPXnRajHcUYHKxi/pwhRBNpSbUcoxJHqETA7Jk1NNodvGj77RDFJey2fG+8/OUv50iQpr5MG17iDR3Eynnwe3dUnm6PKit3zs5CfNmVBec0TXM3kSq7y34YWSOc5/AqLPdsdAZu1MzdqCxqRKogWlDxai8nyJ+S5FSKY2cU4kTpr3trv6qwRfUK9q+CLcKqRVRP2aaDlTjVYNxQXihWpabTwapKOB2sOl4POnR+nqKwP7ItVfAQVk+5QuyiiEGE2EQ0sfKhx6te9WosWrQIv/3NRZg1FGPe7JmoVHs/9xenCarlGPNnD6KRlrD9wnmo1AZx6stfgWOOOQZ8tsZUY1Gj1cOv5TkuV8pdt3yH5Op9qFPQtIQOxZ/zqfLgazk0eDUq99BaZ/BlSB2kClkVWxWCt8J7euIUWosuaoyav6m31UlQqhXC6Iahgn0hWHUcipVC4sqJe383LI0i24pVHYayQuJyrJqqhdK5UO1HsaqCpmmaVd21IOyMg9dNF6s7DDUol6l+3/2cm6g4JwCynZrZ2TjqqKNwwP7748Ybb0Bt/FkgbaJaLqPRaqNarWDn7edg8ewBJJXZOOFlh+DFx70Yc+bMQXfzd7hNnUd35KGxunxdrqH0k6++fUGzA5WrkwC1cc6jO/AoinrPs+CgtFMtSLqw1ct59GSHrJC7slIBuWyrIJKk93secdx9uhSVT6mpKpS2q/3ze90H4hE7hJXjU0G6EXmRUB+Wq5SYbanT4Tx1Op0cVk3d+mFVeqhYlf2pg1dq6wrnzkDP0+s1PdINbU7/Fas/0IdMolKpgKtwnIMQVnXEqsyho4hldP+efI4aRfd9V95Ds2bj5FNOw9rHbsfIxueweNF2+NPqNahWy1ix23ZAu43djjsdg3O6K0pAlK119PqhcwLoMPLj6e8w1FDJQN1hqk3q3PFzyiLE+HzONOipXF0Pyh7tQwqonl8jFRt07wfkUw/Prfy9joFK5hFD29KH8/h5TmtDxUBOvmPVMWkUKMLKf7psWKQAIYEDmIQV6KUonAumYcqG1AGHiprajjpUfq5K4HPDtn0JlFinY7wefIBe7UJZhToyxepBKoqiCbPsHU7daaRFh57Xb7UCACoDMxCnTWzePIwoAirVAcyePx9Ju4OBWfM5AhsT6xPOdiacitmB90sdU11TffEUtkiuyhRch1WumtL6SqUzoglnX86d4AeVT/dDaJ1DI49+74D403n6M4U6Aeqc1MDZtn6W23wkE80x6KaWnsDy96GEsPJ6HYffvcpx6NZZxZqmaRY1yRq0ffarBUpPW1RoWmxyVsNoHcKqBU8VPOcthJWf6RiLsLIdPhy2CGvIGfl8Et9UWPmUrH4sQj+f7Ez4N9Bv3wMAzJi9EKPrqyiVIqRIUa5WUR4YRLk8hCiOgDSZ8DoRfcEUBx1G/jN1cJQj5cp5VFbvhWx95bU6r1pj1AyAc6qMwtPERqOBarWapc+xevoQrSFtBPLLeFqP4HZUXqfPX+TrwMBA5igoPE4KoxcVL5vKiTFwFxn71DsxVRlLpVJGaTUlYlvqeZ3SEas+nZx9h7By/HxgC8fNz6rVai6C+zZbXQ3RcfA+ET2POD2HV6zO1rQ46QZehFXTKDoK/c1XxSrRpi9WVUwdgzp1jXieavFVn8ilUTN/TF72zx/h/Q3Z1RJ9S7UZKJermD9vLmJEmDdnFpB0UJkxa6KZCGkadbkEV1dSdD+bSEGibIwTTiUbYyzsZvLGwmq1mjNuxU1d5BzzUFvQOiB1gTZGXdDVN6+lsZ/BwcGcHpWVfoQe+sqGldLre2UZGsE16oU2UHlu6sbstEmjg1Jcpa+a4wL535rwKKeG6ukTDUmNjc6JWHkQm0d4PacIK9vU6P9CsapDcKz6g9V6OFZ1PBqhnJn5k937YfV6izIoXs+xav1C6zt0mmpUfjjLnMQq8mdPmqve5920IYrLKNdmYnR0FIiABfPnIEoSxHEJqbSW61de01wvk8fK9ESdgqd6QFiuALIal6fhqtuhrMELzpopqL1odsC2s+dZaO7CRjyH5SCVwmhOqysPeoec5tx6HSO0PgPQQVFh+Sg9RlSNflwKoiPTvRD6XguLTv+1JqICYJ6t+aRiBXq30/vn2j7HoVi9fqLsKISVAnV5FWFlf3ovAbGqM+ahzkvlr3rAnz7kmBSD6keob3cQjpVOUA2FuHwFp//RM/4omghSEaO4nZkm6NUa5DVN0Gk3UR8f7xp/p4W4Up3wCKxeyuvE/6Oo13vWrbzneDQgcD6ANChXZZYaANzJ85/OYRdj/icNvYBJuWqQVkaROSjSTKXtNGq+598aadXwtEDJ8wcGBnJK7Pmw5lVUKFdqjbh0Pp5CeFFGBaB5szIc9aaKzbGyfWVRjhXAlFjZJyniVFidDhKrOiFngEVY6ZQ93XHs6uyIVZWGmAcHB3MKqFg1oADI/VQjz+mHlfrQD6sf6kD4PrVNUXpZmq1ShI80nTD2iTlotTtIU6A6MIg06aBVryNiAym6D+5Lk+4/JDaeyf1ybGxAHZTKm/NNOfawdV+LHqIdkiswefOeygTo/vaL6pLWIPl5rIUpFSIb0hRElUkLLaowFD6vU2/W7+DOwNBqBaMOlZj/1HDVE6vi83oqnUatvFfv0fJQfveXwsrzi7AqfSzCqo67CKsqkdcspoOV5zhudTz9sCqTULrsjplYWa9SrByDMxI1SKfwNgpwR2XREeXqCQBrD512HSmATpIijiaMN0lRqpQ0iUEUxUBU6lGICZairKLnFGDj1xQCSJIek1D2RnwewNW5KgtRhqvzyEPlymtUx7V2pfaU3Ruiqw70KEmSZMVKMpAMvii3Uh59QjONW7d9h6JDKHpoBGKRTxWDORuVTBVXdxnqJKuXZTqg3lwflKM41fi0mEis7GM6WLU/HorVi4GKle2HsOo49NDfiGBfjlWNz9MQGqk/cYkKNhVWN+JQbUvHH0VRtprUarVyWEN9hI68QeY9RbcPbUvZCHUkAdIUrVYbnSRFMnFdpVZFHJckn2CbdDrxxL9I2us5K2dB6jTSNL906nL1a5Uxql3oYoEzNM6/snFNXUJyVXnF7snUs1P5WOGngNVoeL1HeJ6rUULpsle9tX0eHJPfg6BjYjVeaX2z2czO9/SiCCvPZ4qgWMmmiFVzaaX9RVg5H+xXV5f8u35Y4zjOsLJtYtU6kgpeV2k0GilWKhcw+VfcPcK7DihWNQjF6gxOsVIu6ph4TbVazT1PgUc/p6FGFf4+yaUCaY5VJJnXSDFRAyuVukyjkyBJOkDaQd4BpfJPuYI5KzqhrCbCz+QV6SQdLpKr2g+AvnKl3N3W9Xz2pcFM5Qqgu4PT6YxHJzVuzfc1+mjlWg3EOyeDyQYwEfmcGmkeph5Q29P1YTXiot/7UCULYfXovK1YeZ6OR3GFsOprCKs6pulgJcty4/K0xbFqcZt/q2LROfhc6ni0AKdYVWY6Z/ycKyBeG1LWqzpRdCjb9c8jFiYRoWu0MSYZ/cSSaPeUDraMbEWnkyCOIjSaTSStGJ3mGLoP2eo6HUTcZ8HKZooIUc8J5ZxXr8904jx1FEBvjv33PlSu/Kf3h6h+MBDStkNyVR0Open6GfUmZsN+qIIAyHkjDlQjBT/P8ps4/4Qf9YRKt50esR2mHox4pKYe4TXPddqrRT6NsK5UnmIoVuKYDlYK1x9NxjEWYeV3pI6Klf9ChhTCqjeO6bwrHo9SmSrLuBSrF5R1iU2x0rmqXHVeOU7iIFa9RgOKMjOVlQYiHuH3aqhME2Df5Vc0ul4lRtJu4k/Pru3qAlKMjzdQrlZlFQS5a9I0RaSrMFm3KXp+I83SjclurxcwPC2l8w3VkHRe1Ikrk/Pgwc9DcuV5+mQ46kXsnomNqPA80quX0kIZ3/Na/hwdD/VUXApV6s2/ldJ7QVInhpOooJ1NuIERq06EKq9jZX/TwcpzGW35yk1LSgcVK/FMhVWXKpUp6Fj8uYuUr2LVZ4U6OyrCqs5FsWpBtdPp7eRUxupzokqtmByrOmDVRZVNZmrBNMXrBZ4+yOoHScfE0WnX0WhP9A1grNFGqVJD2h7vpjIT7ff6iHL/0qyPbg0DEvUnBglEQBpF+VEJVr23pkiuipeF5FCpQGUJTH40X5IkWZCi7Dywx0oz3BFw8EqJVPAUqn5HJWMbIe/H5UMVuCqsGgsVSwuw/Nwdmj8Tgg5D6VuIWVBhtwUro6hi9UMptvapjsuxqlCnwgr0nDyxaiGyCKvuT+mHVdstwqpRaiqsuWJZAVZPmYA8e2Gur05D+0TqxcPJR7foGOWukW+BNEG7MY758xd1xwxgZMsokk4CRCmSVqO7ZNptbGLcAHd+Z8upRduyWK/gv4kjQprbMasO1ovpIWfJudQ6kTMUTacpV2XWnsKx7ziOuz8FoFtpKQAdrN7go/knkE8rPFryeyB/J6TmzipYzYfZ9+b1z+He++7HyJYxzJg9D4ccdjjmDQ1kQLSuEEURmvVRPHjffXh27XqkcRm77bU/9tltp2y8+qPPxKOrBaNbNuHZtcNYtstOk7B2Oh2MbHge9z/4MDaNbEVtxiwcdMihWDhnZm4uOBa2rx5809rV6NTmYd5QbXJK0G7i5msvx0NrWnjn21432dFGEZ5f/RQeeuQxbBregtnztsMBBx6IebMGszlWXJoq8rM1Tz+J2rztMXdmDePj46hWq3jq4T/gVxddip0PPA5/c+px3cgp8mk1xvHoyofwp9XPoZ1GWLrbXthn+S4ol+K+WNkG5arncr60/qJzoVFQI2Q6yQD1tvAJepBOlBDs1HSSU+A18ncEpEkbYyMbcPNtdwBpF8/GjZuweXgL1q3fgIN3GkOp2p3zbJNWxjA0nem/LyT/RZetaK1IA5jKgw5f21I2QbnqwXa7Q+uOSxmmBntlFRzzRHAp54xXBxnKldwr8Tou5QCYFLGcOmkdQNsql8totxp4+I934sILLsCVV12Dhx7/E2qDgyiXSmjWx7HjASfjxsvPQQVJ5vU3r1uNyy/5DX57yWW48ZY70UgiDAzUkHbaGKt38Mur78KJB+zQHQ+AVSv/iOtv+wMOOual2H/3F/UmpDmKz3/svTj78lVY9cTtGCrFaLcaePSBP+CC88/HFVdejQcefQrVgUFUyiU0G3UsXH4c7vz9uaig61ia9VHcesO1eGp9A6969SsxZ0Ytw/r0Q7fjzae/DXu+7O/wg//8aHdekjaeXHk/fn3hBfj5L8/FE6vXg/CSyQAAIABJREFUY2jhbnjNm16H7WoRmo0x3H/3bbjowotw1TW/wyOrnsXA4AyUSzEa4+PY7yVvwhXnfg3gPojGKK658nJsbA3ida8+FZWol+M+etc1+Ju3vBsvP+OL+D8ffyvKJeBHXzsTn/vid4ByGfXa5TjlpddjViXCxrWrcfVlv8XFl1yKG26+HWOtFIODA0g7HYzVW/if86/Dq4/dI5s7pbouV6/5aM2FB3VPHYtu1uvKbnLhMmB1UMONuo2HT8veRhNFyRRRCrTqw1j91FNY9eyG7rIpUow2EtSG5qL+7DBaY8OozFwoDsFrI+FhpXbj2MTur9xJvhqmNqbGrmkugw7no1ar5QqiandsTzdp6RP+vVCtJKCsvzXhtJUdsYFms5lb7nL24A8MBfJVdlUap8dxHOG6i3+Or3zjLNxy94NYsmxvnPaKN+PME47HbjvviGrcwafedzpWDc5GpRQjShKsvOdGfPfs7+PXl12NOgZx3IkvxRe++l4ccuC+mDdnFm675By899PfwOBg18uODa/F2V/9Er5y9k8wWm/hpLf/A37x5c8gjmPUR9bhkx98F35yyc3Y+/g3oNwax5W/Ph9nfff7uPGO+7D9znvi1NP+Bp/74vFYtvOOGKxE+N8ffDvubczq/oZEmuLxB+7AmZ/+NK645V4kaYyhZfvjNUfsgTRN8dg91+H0t70HTz43jNOPOBzjWzbhFz/6AS6+9FLcdtcfMX/H5Xjt6WfgyVsuxKPpHpgb13H+T3+M73/vh7j9j49i2T4rcOrfvAtfOPZoLNt5R5TTBt7/plchnjULUQqkaYL7b/s9PveZf8SN9zyKFGXseuhKHLHTbCRJgj9cdyHe8XcfxXPDLRx22MGob16Pf/+nj+Ls867H+z7yCfzu52dhu6NeitHnH8d/fe0r+OUFv8WWdgUvfslJ+OcvfRMHH7AvFs6bgwduuABv/eAXMGfOEKIoQmN0GKtXr8auy/fOKTmVTWsalLemJV5M9mhJXenqGHdKRghYndhqfgEzSntFxix7yFxElL8UQNKqY2D2Qhx6+OG47rrrgQgY2TqGcjnCdvPmAWk7xxwyRtEjJ1mDQXaTJjq47G2aImeg6lC9+OsMXlkZ09F6vZ67eVPTZ867FqtVBmr/lEFZ8xUVDAejFIiOIhQVVOBKL333nt4nkmMynQZ+/IMfYGjpCvz8zK/gqIP3xUC1kvV1+6Xn4Ko7HsenvvRx/PCbX8aFF16Aux54DAsWL8NHz/wyXvuKv8J282ZP6FCK9vhGnHXW93HIy16DrY9ej4/810W47KprMdqq4u1vew9+fs538dKXnIQk6WDtqgfx9+97L25/6GkAMd7+tjfjgrP/C5/816/jgGNPw88u+hKOOXR/VMu9vPqP156LS256CB/9whn40be/gosuvAB33v8o5i/eG295zSn49S1P4ci9dwHSBNdc8AN88ONnYmujjZmL98Iph+yAj7zzTfj1TffhlNe8Gd//5Bdw3BErUGqsx4k/+QqGdtsBp51wLO57/DmceOobcNGXzsbB+y7HYK13N++1534Ddz4xgn/76NE4+2tfxPnnn4/7HnkaS3Y9DK89eSFuerqK/bYfQpq08etzvoZ/+NyX0EwSbL/HUThwcQvveMMrcf1Da/H1H52P1dd+G/ev3oLj1j6AF7/4BKS1hfjQp/4Nb3zNK7B4wRzEzHk7Y/j7r38bex97Ctqr78THvvO/cdlVv8PLTn0Vvv71r2VzoykHFdRrCxosaAi6GsXCtQainLVnz+wXhxFFZq3KRrpLpqn83Sts5i26Nb4ZC7dfikXPNzFjcADNRh3DW0ZRrdYwY3AAneZW6SSRYdgui5wzo+eQtDA3/u55xO4rUc4sAGQ1Ii1+qjNmKuLX0fa0eOn2qpkFrysr7WOjWhFVGqKOpDsXk+9SVArJwfMzL5QpNUVUw//86rLcWDJP2G7j4vPPQzNp418+9n7suHQZjjvxpfjIP30ZRx9+EGpljq8bdeI4xlN3XYs7nlgPPPFTvPfmS3HwYUfhY//0n3jFaafgN9/8FAZ3OgivPWkFLjv3e/jUZ/8Nc5YfiU988ET8y9d+gl99/TO475Fn8Pef+S984v1vRLU8+TF0v73gPDQ6bfz7Jz+IJUt3xYtfchI+9Nn/xFEH7IxXnnAsXv3Wz2JmawPO/Ohn8d1zr8Dr3/e/sP72n+PO1S289tSXIZ29M3556e9x3Irdszl96JYb8eiaLYg334bTXvNGfPHs92PFnjtnc5VFnQi4+MKL0GqN4pNnvBMv2mV3vPTkv8an/+NUHLrHfBx1yFF46z+djfq6VTjzzH/Ezy69BWd88l9w/Y+/jLXNdfjr016OoZ1W4MLLfo7D990Zn/7ZGtRqNbTSKj71r/+Nk192EnbcbuKR9EmC9oQc1j90C254aA3w0EV4z93XYsWhR+D/+8d/xytOfdkkquvy9YCklFhviFKl1q3lWmcCDTGaYBhIu5ZH1jFhm9lW7mzpkimDpArZ6d3v0rSD1vhW1GZsN7Hq0x3T6GgdADA4GKExsg6z1Ojl/9CqSs6B5OtkwcNSNU81aNQM3L6BUVNAZSDenmYRfO+PgdD+KJOybvphpZT5jl/gS1mei6r3023J7tk0p/W8i9VcVZ5ypYL3fuLz2P0lD2D/FYdgj913xcyBbp6ldzbGce9RbrscdjLO+vpXMLjgRTjk4AOxaP5cxHGEpL4B5//2d1i8+ECc8aZX4Pd3Pow3/93HceYnPoANK2/G72+9D7O3X4Z//u/v4cgDlnfjkWDl2N/ygU9jyaGvxN4HHIQ9d98Vc4ZmII5j/PG6X+Ch1Vuw7Kk/4KQT/h3DmIv/852f4Q2nHoNffGsYw1fehcNf8g68951vxXZzZuSibnXmfLzure/G+z/wQRywvPv7E26ExPqhz/0HDn7l41hxyGFYvmxnDNa6u0Kv+9XX8Hyrhmf+cAVO+PcPIZ2zFN/52UX46+MPxJc3PIjr7n0ax7/7DPztm1+LeUMD6HQ6+Kev/gwf3trEou0WAGkeq8p3/p5H4Vtf+U8MLtwZhx6yAosXzu9uP5JopkVJD0S67wbI17aoH+pIdJm53W5PmOGEwSvXzz6bWKZMLcanasKM7jGTiC7HSLtOpdOqo1mvY87CuYijCPVGEzEiNJstNJpt3HLHAzhg310wv9VAXK7KGNTos//pBzkn4ex8YgIyI/fitqd3XPnTgj3rhl605zyqXNUOgd5Df6mPvt0AQPdHhvbaa6/cmOl1kiTJVVXZgN9mrQJWJVHF8LyVhq5FGM2rtDLL6wmGEYfnaVVXHRpf+a9UKiFK6vjkGe/AVXc9iUOPOQHvP+MMrNhjp0lYOd7pYOVY0jTFmkdvx9ve9WE0ynNw6qtej79/799i3lAth5XCADBtrOzDH5/vWB+580q864OfQXXuDnjdm96Gd77ldRiq5TfQMZJo1OYYVH5FWHMrOFPINU1TXH311dl4d9ppJyxbtmxSoPBVLf2b165ftxbtttyjFEXgRqtcIZPzkRUR8kuU3Qv0yea9ukNzyzqsW3UfluxzHM754Q9x2+13oD46ijSO8ZkPvBbb7bQvHr3jWhx8yuko1WZj8pFI/3IUsYns6xTVWg3z5y+cJFfKiCmKBl3Ojf4UhTIMnueLFypXZ3TsT8sLK1eu7C6daq6jglKqoxFC9+tr6kEFcLCqRFrt5a+x6z4H3zClE6KMhudoBdfplU5ANsHxAL74P7/Ef4jnDmFlX4pV+y7CumSPI3DV9bfkmJpj1RQvVAgswqrFZs/1iXHPw07Gjbf+1aSCoiqC58RaJ1DHUIRV5QP0Ho7EMTlWrT3omLx/bT9Exc38gLR7D0cUxTn2oPE6gkTS7DOg91g8LS2kqI9uQqkyE4hi1Ot1lEoxUkRodxJs2TqOHasVLFk4hE5jFKXqEAHlx6QMQvvUcckc8G++qlxVfhpMQvLlXOodzWTqDEb6aES274fKBOjtBYrVYEhhNMrzUK+v0cAr33po8YRg1aOpESZJkqNOHKQeyhI0tWE/dBweBXVTVhFWVWbP54gztFmsCCvP74fVjUbbU6w+946VyqJsS7HqjzUpG/BakzJCnfsirPp8UjdsVXp1iqp8RVg1EipWIEY6sWLQM8JuWpE92o7/pyMQ/emtXwgDsX/1LRuRpDGQpoijCFu2jHYxAminMeJSjDQtobF1Y7dfbsDKnmmBnPOI2I8dHGOUO7cXkDQ9VXmoU9bHS1IunuprAGCtQ9mhswnVTfabBRYdRCi6OuXVmoQrH79X5+F003NR/gN6G6ZC1EjZj77n5Oot19qXUlnduBJiTTnBRVEhVs3PdX76YaUCKFZnBSGsIcbkt5ezTxqaY2VkUWVTvEVYNWCEsKqDUWagTCRN8w97Vse2rVh79Ybu0f1rokKZ8o7RrtGmSQeTdlFGEwXRyWF+AmMTcRRhxpyFaLVaGB+vY9bQEIAUCVJsHt6KtN3AzIXbA2lbCqO64oJJziEUvemcNCB3V4Tzt5drfcLTUmWInHedZw1StAUNtip3jpNBzuUaRRFiffisVkPZOQWqlESFyIHrvnJVWjV6pbaqIO5geL0v4/iYXBAK3vvV8UyFlUcRVn2+hnp2Xj8drOpQkiQpxBpKIxyX9z8VVj002tOxTBerfu5YncHoeHnP0HSx9tIYoe3Za4ruvRq9/9yp9MBiYtXEagoTf7frW1EfHcHQ/MVodzoYr9fBVYwIQLMNNLeuBaIOksbIxHXaVz6t6P6L82lKeGRZH5qyKXtWOasDD6XbKn+yOH8eLfWO56lcfRWF58RKG0M5jFN50hRtME3T7MYwIF9kKTJmXufeDegpDqO/FsuYqnh+y8jpT+NWOu51gVCE1e8Uq0Y8xUpP7M7Lsarh6HnbilXTEn1+pZ7nhasirDpHxKo/hUesSlkVqzqIflh1bqMoypiOFuv6yZV1EGWVE632Eo80zSh/9zwE3EYKTOzJ9CNNU3Ta40CpgnJ1oCuTUgnDI6NZ8XTG0BDGxhq44aa7Mb5lGNwWn2MH2qaMTY8I+dTL02sWn71WpHJVZs759XSUcmQqqtfqvSaUKw+3Xb6PdTlOlUgFxgijE6vnUoE1D9d0QnMqXkcjA/K3TfN6Go+Oi4qmY+H1OhH8p5SaVNi3tyueflj1NYTV3+tjyhSr4izCyvlwrKoMrmDEqsL2m/z0vbJAb99TG1/P51wzYDhWl6f2rUuDGrlCWNXJpWma5fiZ/sn/VUbZx7nzJs6Z+L9u1+J17foWlCozgChCs9nA2PgYtls4L0s3xsaamDlrCLutOB6rn3kOabuZ63uyM8uPyVO7yUcvleersjm3F287FIz1u35y9bSHxVCVd8w6gUY0rU9oJwQaWuJzmqsK6XSeiqLKr8UVDrhcLuee3K1e0cek7bJ/LWx6eqB53XSwqicPYfVoqz+E1A8rgElYNbdUrI4jhFWVVeWjxqc1JlUspZwqt5Bcgd4+CS45+/wr81TnpMxTH9jrWL2GoduzU9AX5A0vMyB5ddPUJCTTnaSN5vgIKgND2UmNRhObR7ZkTmXT5mEknSZ2220X7LBwJtrN8aADyP4WvQx+HzjU2JVdqNyzSB+Qq/YRkivl5osHOi7KgayS44l1qdIZg2/v1r0Amm9rRNBBh+4F4TlxHKPRaEyqlLNPX1pkezqR7sWdlimFU6Xrh5WfTRdryKloO1NhJa7pYFWh0pA1euvf7kR1vOos2Ycv6SpWb9MdrDqfOM7/Pq1fo6mgOiVtz3UpU+woytUZ0ok9DSF55o40zacjaZq7Lk1TtBtjaDfqGBiaO+HEuitIMwYGgYkb09IUaDebiCKgVKkgaW6dNM+hfyqDYlaBTCdUb12ual8hHfbaEa9l0TJN01x9Uc/V9j1wxnHc28GpnkqVSC/QDjkANuQ3t6jyeLQBujvGeHecKrAqICfE0yT1uqGdZj2dyG991YfXqscMeWXd2NIPKzEqVndijlUrzp5SeP1jOljZRgirKpv3x2MqrHxVrNqnjqPZbGaPPFCsIYPy3Jj9c24nY+2afM5xisz6HblUxBwvADTHR9Bup6gMzkKSdG+arNfrKJcmfj0sTbFldAzNdvf3REqVGpLWaIY71LbOE78LObPQ3Oi1Hqw9XdU0X+da7dkdEM/VVTPtU/tg22XNbXR3oE+CKhvzGVJtIP/gTzcaL8ooJdXv1NGo12s2m5N+B5P9aarhuy31Bhte60JRp6aTzPG/UKw+Z5r7ca51jin4Vqs1abu7pzG6f+PPwUp5qKPZFqwuJ00b1EjcgRKrykv70/lTrGkSpu+hqO0GPJUzaTe2IOl0UK4MZAGqUorQ6nTwosVzMTg4iObWEcTlGYgioNMpYXzzWgxut+ekvkNj0785ttA1nEN1+OoAvBahMtTt3BrYKVdlzz7PWk/0+UuS7u7mMjstysMJjspEwVKhqUyaAigIduqrETp56r1ClNwr5E6tQgYPYNL3PrlOw0IsCsj/XJ9jDc1faButY/HCMr9XGqmbadRBepu8ziOmYlXMRfNArJxn3YUawkqDnwqr9uVj83YUqwYPnyc9fC6KzgtF/ey7dgOVgVlo1rei06xj5LkncOyKXTGjVsFArYa58+dg8ZIdUY4TjG96EpUZA4jKVfh9adM5Ch0L8sVnZ1+h9HsqufJVHy2hS65aE1HdC8k12+7NiKJ5PY2bBSkKj8swSld5nlMgXxLTc+k1uSXV0xiPfEDPcNW4QmkOrwk5EmLlOY5BU42psPoYldJp5NfUpR9W3Y3qWL0AqZ9NB2tIrpomatriQcKxegRTx6fMkXm0yohyY1rG8/phjaJI7+cMGp8qduh7nzue22nVgaSFoTmz8fT9N2N8bAQzZg5hr733wOaRUTy/diMeumslnrvkJrz6FS9GmnQwvHEj9tpzZyRJG1E8uVjYLzUpPCZOU6epKxbuXKlHIR3Wflk/8lRDHYzart6cyddWq9V9noXmPl63UEXj8pb+YlZIgYHJvw3B7/1+CPbvD7ylk9GdgxpheHiNRJVSVxfIRHRS6cQUKyd+ulh1jL4ioVg5xulipTHpoTk9x6GRw7HqdVoncazsS52Cji2E1SOSjlVTFP4QlCu/YtUdpjpmNZA07RUlQ4fOS+i71K7VczvNUYyNbsVTD6/CmufW4pln12H18+vRbHVQqVaxdsMmpClQjSOs27wFO86fhWuuvAUpIhy+8xjKtVneYfZ2uo4ixMzUUevvf6gR64oVAwzfq7w9wOqtFaqrQM/mNZWJ47hbs9CJbjQaiKIoF3nJAPTpwVQWVU71SKpA6sV0n4NGNRqn0y1NZZSS6vd+sG+OV5dftS3+oHGtVsu+/3OxqsP9c7ByjP69K18RVjcMPhFtYGAgw0psHIs6ROJRBtgPqxZJFav/ktmfg9UNnteFzlWHqroT+r49Poynn1qNG265D4899RxaaYp2miJNI0TRGJIUqERAI0kwsmUUO++4CBubKWaVmug0x7MbyrL207S7cmOMJ3eO4fKDc6hy1Z3Rek69XseMGTOy+VEWqzUf9sUfVVb5eS1Ra38SLOKs2JYkvV++ovA04ig9AnrPrGCEZmHMFUgniTc1qVdTQ9SIr4rrdEzH4ZTPI71GKTVSPrZeU7E4zmPlGHpYI7RbzeyJS4rVqbZjdafTD6vS8ZySm3P0orCOQfvhPo481sk3oTlWBo7pyDWUC3tq4mPthzUUCPRwh6CHMiTOb8R/ZrCt8c3obNmEmY1hxFE6cbdHdosaAKCZpJg7ewilTge1Wg2DM2ZgYKA8sSKy7UVXP89xKZNQJgxM3ovBYAfkFyl06V+/owNXR67nOzvOVizf/e53n7l48eIcFVYlckqiRuTVVZ2AkDGrUioN0pzVB86+2QedQalUwsjGtXh6zQbMnTu7G9XadZz/03NQXbwbFgzVsOaZVdg01sbcWTMRRRE2Pfckfnzuxdhrv/1QSppYuXIlakPzUC13l8cevONa3Hj/auy7xy5dRW418OC9d+HXF16AeM7OeNGi2bjzhivw7bPOxn2rt+Kog/bB2JZNuOfuO3DlFZfj8ssux+9vvBnR0GLssmQhoijCumf/hHXD45gzq/sE8OH1z+CcH/0Sex54CAbKk7FyTupjW/DYY09gYGgOatUygAQ3XXURHlnfwS5LFiJN2nj6iUdw/XW/w6WXXIKrf3cdHnhiDQ48cD+U4wiNsRE8uepPGByahWq5hHariesuOw/PjFax8w4LUS6XMT46gnvuuBnnnXchdlh+EObOrGB86zAeuPduXHn55bj00svx+xtuQnnODthp8fxMvluHN+D2m6/HBRdfheX7HYiZtd7eAHXqdDqrVq3KPps3bx4WLFiQcx4qV9UvMhWeNzY2hiQprtoXsYvsfcipdJqob/oT7n/wCdzxyBo0OimSFEhSbvzq6XK90cLsObNw4D67IinNwi47zkF15hxUZm4HINLsY8rxhI5SuYSZM7ssRYOpOgogn0Y4G/N6hxZI9UfQPZ33MaqtRlGETZs2dVdDNDdSulmv17OBEIAXRrxAkitISe6lHp7FGd0u7A8CJv0KrStHUYQ/rbwL3/reT7G5MYgvfenzKDW34GffPwu3r1yPY05r46ff+xrueuAJLNnnWPyv970Bzz31EL7+jbMwY6eDMbr2cXzzRz/D6jXr8Op3fBQnHLIrbrziQvz8oqtw2uln4N7bfo8/PvwEHnnkMSxZtic2PbcGraSFy391Du56Zhw7bT8fM+bMxLnnnI0/PPQEdt/nQBx8+HH46xdtj6vO+wE2DI+hPjqMay7/Da654Q7MWboCn/nIOzDy/Cp84xvfRH1oNzQ3PIWb/jSMYw47IIc1TVOMbVqNr379LKx5fgPe8/F/xQG7xLjywp/g/CtuwXs+ehhuuOo3uOnWuxHNXIDDDz8cbzz6BNTXP4Ef/vpWpGmCh++9E788/zdYt2EYH/zHf8PyxSmuuOBH+M01d+EDnz4B11x+MZ559lk8+vgz2GO/ffHc6mfRaY3iwp/+Arff9yiW77cCBx1xHF6xZBGuPu8H2DA8irEtm3HP3XfhgQfvx6rVG7HPvnthzeo1aI6NYEtSxZx583L0lbJUpaSstRYUSkl0T0dR5A0Zn+qlpz2hCJ+m3aehtxp1HPuy07D3UX+Fyy75LR54+FG0O3I+etxhy9ZxlMslHH/iS9BctxKdxtaJNifvqdCjCIdeEwW2rpMVEoPWAt2JNBqNbI+LbtDSedRn4obGowscymo6nQ5K73nPe85csGBBbgLZCTvURniOey8dkAtMVxO8aq9LiO491YHp+Lp9x5hZSYG5S7F8uzLOPutstEsDqCcRHrvnVsze5UAsKNdxwFEvweZV9+BHv7wUM2plVKpl3HDjbTj+r07G2mfX4dRTjseVF/wU9zy5Ho0tIyilY/jjo6uxfO/98fo3vhFHHrgbrrj0cqx8+AF0Bpfgna9/KX598aXYPLwFO+yyJ97+znfiyEMOwJLtFyEZX48f/+JitMY346qrr0Nt7hJsP7OEPQ89FummJ3D2Ob/C4OAAypUSbrrxFux10JHYcdHcHNauQy1hwdwhPP7cOE45/gD86pzv4smNTYxvraO+YRWe2gy87k1vwStPPhHLdt4Js4Zm4pqLz8WzG7fijhuvxeNrhnH4iv2xfryCk45Yjl/84Gw8syXBWL2Nrc8+jNXDbex/0OF48+lvwrIFJVx+/e14+L67MXfJXnjv+96NIw89EIsWzgfqG/DjX/wWzbGNuOqa36MTVbDfocfgzW98HRaURvC72+7F/ff+Acv32gfz5szOFE7z4DRN8dRTT2XymzdvHhYtWpTJXwvqqhf+eZIkGB8bzdHsfmmIG506jOz8NEVz61qMrHsGc5bshcU7LsURRx+D5bvthjXPPINNwyOIIiCOIiAFauUI5XIJxxy+DwaGtgM6LXSaW1Cb+6LgioiPIeTc9ChXypgxY2Zma7Qxf0Se2pWmWkwX1dZCfbOe5k5UWZwuoQPoMgstbvBCpS/6+H8OksxDi1ma4yiFouPxDVhUCqXgjDhaW3BHxf7mLNwezz75KDYOR/jW9+/Hy1/7VuyxqIKrrr8Tex14KHZfMoTPf+4yrNtyLsqzFuP9H/4HbH76PqxcPYKj3va3GH/6bmyuN3DWV/8bexxyHD78+mNx/RWXoDJvJxx95KEYrE5E+Y3rsOyAI/HSk0/Gzku2A9IEn/rsP2PO/AWI0vyP5wwMLcBrXvd6zF+yFLsv2wXVUgef/8THsGZLHfdUZuFdH/wHpBtX4c6H/4TDjjgaOy9ZmDlMlUNcGcT4hjVot7biq//9dRx2wsvxhiP3wZWXXoYFS/fEEYcciFKU/+2Hg446AYv3aWOfvffCwvlzcONvfox2fRO+8tVv4/ATTsObDtsDV1x6JbbfbV8ctmJfRBO/u7Kh3sRRx52EU/7qJMybNZhjBpUZc/Hq/1vb2fxKcp11+O3qvrf7jmdsJzbBxMSOgx2DCJDILGKQAIGUBQs2EctICIl/gwUS/w4CCSRW2UUi20iB2IgvoSCRxPb4Yzz3q7tY9DzVT/36VHffiSlpNLerq855n3Pe836cc7rq29+uX3zlK/Wll39peM7nfD6vx1fr+sNv/XH90e//Tr34/IPm3AOTazgElM/zJY4uHNl6EOy8607ZD3nxqcHa+vv28qPq+1mdXdwfnrP1q7/+tfrNr79bH3z4sD5+9GltbtdVbPG+WVdVV48/+O+azxe1ubmsfn1TNT/bKzvToGNpCPflCpxTkUzfuCfbxA681U6ez8rUv2q8fIpMs+9973v9m2++uTcz6k1UuYxFJbZyns/AaFj4qt2255bALiutJue8hbmq6ic//o/6n/cf1xuv/0rdW+0ekz+fz6v6Tf3rj35Y3b3P15e/9MWZMtTCAAAb6UlEQVQ6W4wfT7e+flQ/+OG79cpXvlovPPfMUF9ua+aeu7DOZtuVluVyWf/2Lz+o2/Pn6rVXXq7FfLwOTtkt1qtHD+uH7/xnvfbGm/X5Z++NlAL5/Ig0e9mu6+qTD35SP/r3H9dX3vhqfe7BvdE9XNtipSzPGThNcI6crByegJvP5/Xd7353kO3VV1+t119/fa9tvYPQ7Wy533vvp3V9dTXizWPKi/Ndnv/wv75fn3z8uF7+2h+M6v7Hf/j7+pu//bu6vV1X9dv3nf7e736z1p9+Un/6J9+shx88rNX5vM7nm3r21bdrce9zezK4PY/JW1W1Wl3UCy/+wt5Eca7iuY2rdnMYbisbHcuR/doyKOgQW/dns1m9++6728jCXsCGgoHsJx0hZM4luFHcKVbi1Wq1pxRsb84c18t0DAgeSkqZX3j5tfrCy7uGGIVXNas3fu03npSz/4LY2fJ+vfXWW6P5lJubm1GeZ75c6TiV9bU3vzacZ9s69+USpAfm+b3n6hvf+K3hs8PSPVZ1NJ1/77kX67ff+sJQvo0aS8M5T+V2zP0tT9OvGFjqrqohAkFWwmza2fX482KxGLZ7pxM6dBwyGv3N49rcXtf56tnyNszNZlM//dl79bnnn62HDz/ebsyrqsurq7p/dlYf/ex/66Zf1j99/5/ry7/8oL7+0icjY5H18Pexw1GBo3yz2FnQjl6mdr+2dDj3V7Tai7Hofu37Jw+/aeWM9ua2ZoZwwev1epi8MrgbKZ+61HXd8CAZylssFsOsra/1ZiDK5ME01GOGXF9uMcDKeW9wseXOulusmf+ZlfNYaWSG1StBDj/dD6ewHvI+yJ+sDmdhtQ7AiqFusbLr1P1Nv+LlmJfx7PwUK3W6vC3TaWnH1DFqn76vm6uPanN7U+fPPF9V4ur7Wp6f1c31bfX9pmbbKYt69sGDevbBg9rMzuulV1+vP/nOX9Sn7z+sm08f7rWJ63ObTaUF2+v35bRRzekCf5cRemtlqmo8n+F+TTnRU+qbz+e7B/ZygoJt1b1Mg6B+1Nx8Ph/mGmwV7Q2t3EQrXNPahQmwJzfzfxTSnsgNdH5+PpoTsSyU67kRsxPlYDA5pliRq8XqtnTOyfeUa9ZUOFimWL0sZlZPHDMTnqzIlaErE9xd1+0tbZs1Fdvt5xTGnnOKdTabjfa/cH69Xo+2M7QGYGvATn3XV9XNow/q4/d+Vsv7zw/X4pg+/uSTqlnV7Xr3WL3333+/5ot53d6ua9ava7la1Zdf+2JdfvLRngGYSjss1558Zn1yoGtVY11yvxKtUaejPDt99yvj1ikxhx2ybcACy2IL4heX4O1zUCGcJ6MsuCvMFQ/nYQBbwe1B/VhzzuVvGByZEJHkfhEUIbewetsz90+xZqg9xeq3O6Uxm2JlcLneqvG+frNW7VLB/GUiCmIDb1baYWqugDocraRnItU4Pz9vRn3J6gGSs/Quz33oMHqxWFTNqvpNXzzYdihbA611tCORvm6vPq5+vtxObtrA99sH7Txz76I+/fRx3VzfVF9V9+/fr9XFqq4vr2qz2bbHcy+9Ut3Z+LcYmSa16resw/V91Xp9W4vF2eDV3aaeu3BUZp2nXzOqdL864s00hRQ1+3U2m+1+derNGg55MkR1RIDArfVcd7Sf2u2UgjJct8NZGiJzWb/s1YaDMqg/O8ShmjvxVFZkys5OVphywLnuQ6yOQPwyoFYoyeeWlz/EaoOckV6L1UaP8s/Pz09mtTF1me4zszoKGaLP0asIt8/S3A6yvsYvRO5rf3xuzw3l317X5uaqLp59obr52XANZWw26/rwo0d1dX1b89l2D8T69rZWy1XdXH1Y1W9qs76ts4sHdXP5sPrNbdVs8aSMXTkpz1TkyP9dNx85A/cJRsDphvWddnKb+7dZblfqdLpPGa1+rapa5A+9PKHpQj3Y7P18v71pLgc6CrEi+MlTDHAGKvdkPuwoxgaKa5z/WsGp0/IkqwdFsjp0PsSKHP671aaewE2DZVbSJXvrZHUkaHm9qpXzBU/LypHG4RCrDbWjuxary/U1n3/hxbpdr4dNUlue3Zu6bm9va97Na71hrooyNsOGp03fV//kVQEvvPCtWm+qlhfbN5fO4ZtVfefP/rzW63VdP3mqVNd19eD+/bp/76JqfV3nFxfVLVbVvfRS3Vx9Wuf3nq/tk7xrxLB9AVL/5OfnXa3Xt4NsXTer9XpTXbczFO7XVgRG+3oDXKbDjsTdr3bMzCflfFGOMTvQhQeOC80w2bP1OdNtQXYWcgzLOe/hQClZ07XXQVDnaX4YiBspvaHTkFa5VmKX70GPnPmcBSu9WbOh+ecBSYjnNM9yfNasNgw2EBw/D6uNE+ddl/v17bffHup0KkT7tFjtWAa5F4vhtx02+shxdrb1iIt+nPZ5Tgz5tu30zN4E4eJJdPP6G18dZLCsHiuDt3/muVGEvR3QZ3t6sR2YF6Mfci2X43HiCJx6HEm6T5ymWDY7gpw/ch9yTzo5p2Sj+RJbH1/k0McDyd7BnsoDY9w4u/DIoa/rtQXLRvP3WFU/tTvDOA57axu21qBusdqQnMLqc63VAed/bofWgDSrZ6TvwmqDkAOdeywXrPAeY/X9GTF6cK7X2x9enZ+f12q1Gu5N5SYK8iBpsXrOKx1Wrgg5TWvpVqtfnTq5fU9h9XfIYxmdQtyVlb/pj/whoI0E8tuwwevoMdPAqX6Vju08gqMAjmy0vH42201MWVgPmPRWrY7j4Ht+sYnwNL4fRpOTP9nI1IOcGZ4dYnXnuAy/AmCK1Z2YrK3ojV9smpVlLQ+uQ6wpp2e5rTjIYyV1GXyPDNlHVqK7sPr+HNQsQ7dYW84n5WylU/aueS7LqKoRqweMI5vWvI1ZKa/Fyr+nZfWgp90899caw9SRTtHL0i3j4PFjQzc83TtzZl/I34S8GSYiON+7E9ypPp+GIxWYcDX3SvA3A8yKnBN/9j7ep3BXVofDlHuIlTJarOblGj87hOtQpCnW9Pb2YslKtGPFslwoUMurUkeyJl8qqY9R3quNZMdYKdd9cBfW9NpmzRTFrJ5Hcz+Z1Z/NPcVqI07dyH6I1VEQ19sgeeDb+FMezjUjL/TtEGvqfecPtsYedPm9K6Wz04Jx2BM73Mk8ifOezeX/6+vrvcnM1qqCZcRQ5DMlzOKOP8Tqsh1dpVV3hOXUwaxug2QlcnKdLVbXiYKiTPaMrjMjE8uUDsBlmhW5GVBuPw8G1+N2dDvDamVN1jSqyepozP3XYk1DY9laKY2P3HyXcwnHWBmU6KJ1KfvVuul+ahlzOw9fb1Y7Rs8JoZfpxHIz3MhBsenDjWyF5n8PDpSIRlmvd2/o4p+fych1GJWpiKAFbSh3Vl5Pp/rzZrPZe8CHWd3wZvWgwKozgKdYHWHB6jkHs6ZST7ESvbTaBsOUUZRTLdq1lZL5vOtvsbpd7C3t5VpPIzvESr12Tndldapl1vSI6XWnWNNI50/DKT8naR3xTrG6b2C17nG9dZh60cFD/WpjaVbKx8BmNGbWdHSwEhwsyKG8pDKbzUYztj7vyAIIGs57HuhQBo6tp58X6Ws4AM6wLr28O8kyWlHyM1zHWPnfuaI9EuGdWV0f13Hez3CwzNyTrJYl89Xs3LuwXl9fj5zCKaxeYuMeO4+nYbWHTlZfdworXPl2Pc4xODnvup2f06+eMD7G6ujmLqy0b4vVfPyNfMmF/PR1i5V/XEv/m5Wys629tN/5cWv2tlZ+BOVmX5fewFYtFYxGsrXOFKLl6W083LmegLJltTXPMrxpCoZWOHaI1Q1P+TZUGUU4wjqF1e3Hd8dYLQuHWbnWSnSM1R4mvdRdWN3PGeK3WB05HmJ1+d5I5D7KFIZ/ZrWnz8GTrJzLe6dYk9esjiDMCq9ZzQBrftdizb0wU6z0YSvq5N7Oymeg/GyDkJMsHshpzSycUxdbMf4RWhKOudHS6zLwsXz52wV7T593Lsx1bqC7sLbKY97ArHSElWSKNT1oi9XvBM0OdWiceX8ac9dlea0oU6yEs6ew8hsTQuFU/hZrGvcWK+dxSMdYqRd5ne6mIbD+En0i311YLWcrcrwLK3JmGn6ItZX2T7E67XMkNIwVey4rjy9qWS4Ebd1btQ2BvfTnjvK9Fta5FE/ATk+aFi9/28F3lMeRVtchr1MkDzaXyeFVAQ8aHu/vbdPZOcdYs3wroVk9L5CsGbK2WB2leLCZlUExxdr3/egtcaew9v12KzGy5jJ0huNW4EOsVuwclBkN+jrX7UlJGwVYeflzi9WGhbSee5DFcxEtVpeNTI5a7ADMeFdWGzvrOxPORC4teYYdnDkhaQXzBGQqHvmtDUVV1XK5HAlng2FFd9iWoaytdVpLg9LZ5IE0VGunJJ1DJ5C3ORc1q7ncTh5chIWwZvjrzj/EynmHl77vGKs9NPclq5lyYtkDj3uPsSLTFCvlULaV17+oPMbqPnH0Rzhtec2a19ggeqAkq+W24Wyx2th4vsOsjkDSGHA+x8kU62azOchqGc2KnPmOmWR1+jn6Pz2Rw07CKUcYbrTWvdm4NKAFQHjeUZKD0o3qCIf73HhWLnc+ltINwOGOoO4pVstsBfN8SLLaunOeyCONxNOw0ulmxQP63lNZUWyUMdvMk88Z+bRY8VDkwKkzx1jt9WDlmlyCPMZqZ3ZX1lZEm/rgBQKXc4w19fFUVg/wKdasJ41li9VtnykbbTQ8/MaAtnQOQf2dlcUFp8Hg3vS28/l8eB4F16NofCbMba1R2+PY0LizMjpyozi6SdahcQ6wtoxjtpNZ/YyGQ6wYOXMlq70fDGmQHR6b1V4wvbWVzgff2dvbayYrD/Vx3X4allcoWv1q2c2a3taR1RRrDkzO5/Ijh/v9GCvleMKx7/shDem6bhRVHRr4+TkNHaw2WpYJVk+2nsrK3xkNZRS1yMb3YElr5JsdXtmL8L13yRnOA5YGSkX1cyLdMS6bweVQK6MURzHIlsu43EdolulDshLGTbFa8ZPV+W7f7z9TNFlpiylWpw5mpU6zWpZTWB0WewDmw3ZPZaWdzECZ/j4fDm1WBoRZ7QxarF6ibHnPZMVAtPTwFFbKY57GTsbjqcWKkUpWD2TKod7PgtX7TXyPy9hsNrXwu0yzIy2QFdhhJfmTQ/bcbdb3/ZByMFtsI+Qc1dA5QJHFE2s2AvZeANJIVTvv5nNuoGOs1OP8NFlns93MeUYTnqzKPShmddh8jNWex1yOWtIY2DFYDntR9wMymZWDMDyf5GWlZbLSrG5P+KZYkcuTnk/Lar21waMeG4qMWoiEeBRijpEWq/vIkV2+HHuKle+nWK3PrbY5xOq03e1FvTywd3hiGopNwW4ALFvmYzx8pmo3WeglMWZTnd+uVqvR4KHR/G4SOosDeD88hzAvZ36JbrwJyYrf97vfYGRI1mL1SoWNmFmRzddTjwdPixUGy2cZT2X1Obdba6WCPuEcno3yLR/KjnKmgiPPYrGo5XK5ZxTxXAy8Fmsud0+xdl23F+rb69HnniA0K07KKViL1SsW6CopBf1vVtq3xZo6nEY29cis1gHKmGK1HHY66dTMil5xH20BK/esVqvh+vV6vV0NsWJaaATB2qa1bIVGdLqVwcqTDWgld16e4bDP2yPSQVZ8ZLf1d6h3jBXlQs6MVHLwmTWjJCuUPWbOvnO+xeq0ocVaVU1WD8JTWZ3a2Bu7Hzz/0zK8p7La47VYvVLgVM+65nC563Zbw1v99DSs+QSx1GE7JctvHaZ+n8f4UoZZM7qjPvddstoQJ6t1ocWK4bAONVdmKIDOcEjiAi2ULTaAgNFoGAyEdgPbCFC/G8JQgOHh8Yie1PFSkFOHVEiun2J1vuhGS1ZfX1WjTSxuA4eEyORlz0OsGFcMQ0ZyZuXeZO373ZbeTIFarJkSwpusHggtQ4pMZs2oosVKPTYKlHOMtWr7qgU7HOSZYqX/7cg893AKK3JMsVq/T2VNB0l9LnuKFd5DrE7H+N+slsd62hFm+lFohs1cBnAaKicouZ59FjSAc//sGBrZZbiTGeC2knSSw1LfQ71WUFvQFiufk9W5e4t1tVoNZRxixfM4hExWBrj57JGGjot78peRKBveywZ/itUhuY2Lrzerr2v1az7+zdGi5cYgc51ZW/3aYt1sNqNNUL5+ihUnk3Nd1H2M1W3qHbbZ3vztn99nFH0qKwadB+qeyprpxymslqfv++pyHiG9on9E5NDGu+i8bMigzrAxQ9c8mCjjHpSG+x09eI6B65HBymILSkd+lqzIciqrPZOfM+AB4pzVA8lGyl4nozdHTDl4aVfaywOX+83qtqTNvUKQrPZ8ZuXHa+7XrBcjm2mc+/X/i9XXWieOsbpfke/q6qrJWlWj5XGvlnC9dywnK3JlNELZjnDMisy0Y7bHIVYbndlstnuehWe7HdoxWZkPycjwjMNPaEZABHG458P1WWCXY0WkTp6HgNw0DJ3Ctc4p8e5eAjzESke0WL2z9BTW9CRm5xy/J0B2s6JkNnrInKwc9GvL6zu0RxazenCYFcVMVnu31BEOs9KvPt913dAGpFDIAavleFpW6qfOvfxcA97RxyFW6xL12+glK9EGBtU6wwupHHX4b1izXWFNQ5WsltdOa4q1qnZzFjnRkpD2AE5D3GkO/VuW0ILkvbmqYEBbR3ssoiKWdyjr+vp6z2O7MSinFZ20WB0eJyvln8patTOoOeGFYk+xEnXclTXlc6iZk6Vm9QrGqawOf630lo/vXLe9HO1j1q7rBtZW+O35FkcnLVaMnCcjzerxYFbKzvQWo7FcLpv9amObKyWcPz8/H014suPXrNm+U32RE8OOklusU/3q8VxV23edZv7kEMuFVu1CP/7mGiBt6anQ5zMvzWWrqQ7qut3ymev033B48si5f3p0c1n5bIUdslGeWdPDtFg5mGjM0Jm2PMbqgQurQ3I61yGkIyq3F/+3WCmvxZoR3hQr0RtKb1aXZVYPRg/0u7D6PntWs+ZmOLMim8t0Gb7e7C1WRxqtfnWq/Vmxpg77t0HuJxsU96sZkV9jv9uzXu5Qw1pQr5G7IoNgNW2Nbf3trR2CAUt41ve7ST/fg+wt7+kOsiJThg+z2lPwHee5n/MtVkccLVaMWYuVGelTWS27lcN82bfZr2Z1lJWsVjanJM6zPehspJN1vV6PWD0PRfs49TyFFS/q6+xwYM3w+xCr+xVW61XKnaw4QadV3NNqs1NY0bncYJis5nV7IH/qQLL6TYVDioNwhGlpTQBwI9iiOi3xbDBlOuTme3b8OQVx2JeTNEQgae2xwDZatrZubDeiUw3uc4Q1ytO63fKhQ3XmDsxqg4EBZLs28riNk9XRVovVKyiZDnl51EpAm3DeslkRXNchVurzVuVTWTM9MKs9tVn5zP8t1rzOg54dl/akU6zWYacvzt2tw/6l7xSrdcTRo2V3fx1jzeus17ASNbWio5xGsLx2rtRvozj6IZnDVneW8x0roUN+WzwE8BKlO9HPoPB5W/2pweoVjvRiuSJieFvVZDFDsvoeK3bXdaPJNORqsWbnflasdL6VICcifUwZWofryUq5hzZFncLqz4dYPVCRHy+arJ5Mn2Kl7Vqs6Ev2q9Mx606yut4pVkccU6xEW1U12jFrZ3cqKw56ijUNhVOUNKZm7bpuuxriLc0czhuvrq5GAyoHXzZ85pzp3R1OOTTMiMKyeKXGIB4c9tZuAB+5r98dU1V1eXk56dnNau/MYQU3q6MAD/YWK6Hrz8uKMZhinc1m9fjx473BkOXaw2R60+pHRwhuL7fJMdaqOonVBn0+n++tgh1j9WA1q70/8pst9dWMrbTvGKsNgXc9w+d7GGNTrF3X7bG6jDTC2SfJSrtsNpvtMzizYTIctLAOX+1FOJ9vPc8KKd8DksZ0NJPhsweVO8rGi0b3OnFrMFNHsuKtHELa+8PLebbbplJTV4sVmTLMbqV5h1gZTFOsNsJm9eScU0HLnm1SVXusnhRvRZpOAzPqarHC58EKY4vVhsKDF1bqoU2Wy+Ugk+93aE/ZLVbK8UDOiIR+bR1TrOiKGYlCUu/M7HtbrK30O+coYHWfT7HOZrPtDs6smJuzAa6urkYhvhseT5ae3NBuyOwsK7EtOHKkR2hNTnmLuRvIE1CHWB2mXV5ejq5ND4ri+uBeG5pjrL4GOZDpEKsjllNYW16mxerw1awZoXAv/2wkzWElPsSKXL7P8md7uV9aumNW9/Hl5eVInszbSeWmWN3nyWqDnWlAi9Wrdq3oxtdTn9OkTEdcx3w+32MlQnRZOVUwxVpVtUApbXU8sWHFyuU8H24UOnc+nw+79+wt3Hm2ykAgB57JypgTUN5w43owXtmJx1i5ZrlcjuSw8coORI6nYfXAdDTVCunNisc9xJqGy7+JmWLlnFktw11YM3JMI0TZ/o5rPYjMWjV+ZmWmfd51azmQ9VRWdCN1mMldjinD7yjSY8SslEc5/O0BTD9lOb6OzWvpXFer1SgqYRwla1UNKZJ326JXsHVW0AxjPQPufMef3cHOs7xOnJNZHvgOdTxT25IhPTYdZUvruYS00mzqmWLNsNq8LVYa0TPhsNL5zttbrDmRbFZHFHQ0eaaNS7KiQFZCD1ob22T1QOJ615nvqzjEmnKZlT6CISOqKVanHHz2e3GT1bp9F9bNZjN6lYJZLXeLFb5kTf2mf5wOIJONqvuV6NmsdkRmbc21uA5YPSnqaCfHV2cQF2QoviccpZMyJHPj58NZ0rr5OQG2drnswyBqTQzRWc73bDCyfD/ODcXMgWlWz9e0WJ3+JCvyMXgyYoLVcmB47PWPsdrQIZND6awjIys8sFmd9rncqt1svVldZrJSt3Nfs2bIbwfBd+kwXCY6SXu6jmOstKtZGVywZhn2yF7FMGsrYlwsFqNJSe5hQLb61azoNIM5Wa1vZiUqO8RqY8U1yVpV1d3e3l5hAPgSga+vr4cOdWjk0J2DhqATbFQyRAMgI4S8xpY1w02+59d3XOefw3PYkzAYM5Qj/LorK+2VcpnDhsb5cYvVEZo7Cq9uD5msVk7kS9aqGrFage0tOTxgp1htNJLVoXgOIDy5vSLXOe0wq3nTkxMB0Fawom+c8yBJVoxJsnKf29qDzylVK+U6xJrG3vWa1U6pxYpxa/Vr1fjFTzmR6vJarDc3N1eLd99996/m8/lfrlarpcMWXodGnpcKno3OZ2+AybAJWK45Pz+v5XJZjx49GhqXzS485AXrfXFxMSiHwyZbxs1mM8h6dnY2nLPiun7u53VwZrWRsII7FeEdGF6Cy9SAAb5YLGq1WtWjR48GheCxZXhIlogvLi6GtrABpH7O88Oqs7OzYatxRgZObfp+uwwOK7/bgCHD/qdlnc/nde/evXr06NHQj8dY+WzWrtvu77i5uRl+d0FZDEx7QuvEIVbPuVivqW+5XO6xpvPBoUyx5kbDm5ubWq1Wg045JaFNeNcOD7JusXI984fIfnl5ORgIntJGm7P1wW3TYq3aLRIwHp9cf/3OO+/89f8BLhwUw6NH/AkAAAAASUVORK5CYII="}]}
