{"current-slide":2, "aspect-ratio":2, "slides": [{"background-color":"linear-gradient(to bottom, #3689e6 0%, #4d158a 100%)", "background-pattern":"resource:///com/github/philip-scott/spice-up/patterns/black-linen.png" , "items": [ {"x": 385,"y": 750,"w": 715,"h": 220,"type":"text","text": "","text-data": "U3VidGl0bGUg","font": "open sans","color": "#64baff","font-size": 21, "font-style":"light italic", "justification": 1 }, {"x": 89,"y": 439,"w": 1322,"h": 403,"type":"text","text": "","text-data": "QW1hemluZyBIaXBzdGVy","font": "open sans","color": "#f4f4f4","font-size": 28, "font-style":"regular", "justification": 1 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nGS9Tcxt23IdNGrOtfd3zn3PzyTGJCgOsYIiO0BibH7yK5lEAhwCmCA6oREEQiDRSB8aoDSQSAeRnhMadBKJBghEAxABJJAiRRD+GjSiBGggbIgITuT37vm+vdasojHGqLmOfS3r3XvO9+291pw1q0aNGlUzfuPf/0/9oe/88G/4k/P5zY9hHoGqqrwiYqDWQswDQBXGRK0zYj6Q5wtAAQACgRijMCby+hgjjsQIIKLy/BjjeCtEALmAMSvGQK0zkIk43rJqDWQBY1Rd14gx+MEoVEQFAqgMflkgxqxaV2ReGMezkPvv+FuoiDlqnYkIBCLiOKqqUNcLcbwBuaJQFTGACFQuxJiodaFyxZgHqqpiHkAmcp0x9PmZq2IcCERUoAKjEIhCIXJFxagYB1ArMhciRkUhClkxJqoKMUZUZkREVVXFmEDy50cEshIxHxW59G4DMR9Vlfy5dWE83oC1UCNqzAOVK1B8fT7oQjy+qbreIysxxlGZF2JMfqTXABEYB1DJLR2jUKnnnAEUEKMqF6IQGIFcV4x5JMYMVHFvI4DS1o1ZqNKf5eBzAxiRQZNBXmeM+ajMK8Y4qjKjUBjzAQBVlRFBu/I7xxi0tdJOI1BrxXi+Va4zAijEiKqFiMF34IchIgoxgKrw7+b1AcTAmA/kOjHGrEIFEogRhQjkujDGBMbk+2UiHs+sdQ3kBcyjwG8JZAJjVl7nGPNIZAbm4AMUwmcGY/JMrYt7dTyr8hqRyXOGqhhH1PmKmDNRFZgHAlGZF1CF0FlFJfRe/F8kap2ImFEAbctnMSYQwLpetMt5IAD+XAwggFwXAkDMR7/T9f4r/+fHD/6/f+345nt/27/19uO//3ec54n5+Iy83vcCI+wsUFXAOhGPT8DrW0TQTqoWEBPj8Ql4/QA43mTfB/DxK6jjE2IcKBlqRQCZqPVCPD6hrhNAIuYb6vV9xOMzcp3gi0RvasSggcwncr14sHlIYCOLmKi8vCU0gusD4/gEVKGuL8DxSb4oaTLjAPLiBq4LtU7kPBDjsT8rT6wCxvFAnR/AOJC1MOYTNSZiDNT1QlViHG+oSn7F+a73efH554PfW0CtDz5LLhQdKO1HBy8en5B5QQaIGA8gL653JWo+efCrkJXow0nnyjU53vgO5wfq8WaHDVQiq/h5CMTku9IpHfS41ws1xjacAnJ9YMw3YL1QNEKGizHpcOV8g4EDEfyuygsREzEn8nphHG/A+Q4cb4hatC0AUQXMo/cn5rPXctgRIfmOMfif60R8+h7i9S3PLAaiEj4FgOyYhxC1Lu45Cji/IMah9Uvtx8W/GwcQE7FeyFy0bwQqT8R8ArVQmYpRDDgKTlwf/Qxi9vogF6oWYj4REcjzHVWF8XhDXR+0x/ngM60TyAvx/A7PZBzAPFCvb/l5Y/Ze0zEu2mwt7l0M/vkYsv0PZAzE8QTOd67rOFARPJ/a+3r/FWA+tOeFygsP5K+LX/qf/uQRY/7m8/0LqgoL0T9Q6+SD2/hqAQisjy/9RXz5Qjwm8jpRyVjVXj+LBlDcJBQQxxuqFnIl4iHjxtRnPoE4tMs8XHW9+uDCWGY8+ffjAHDSNWYBA1xUeVh+1sVFyQXEgYiJ9s7j4N9dJ+J4oK6Lnx8Hn8vvCDkqDH3m0ME7tF76Ox5RGbNgTiad/zGRme2IK2s/gxxIQIctQp/n/z4Q8ymjBioXxvNtO9HxoPNeFzd8XajrAzj4vDGW1gUAJoiMgAw6SIwDWHQkfHcAR+ighg5HoSpRMXQAHorYimpVKMIHgZshJ8CAWihgJfc6+f4p56zoh1oXRkyu47qQAkl2GL2o9BK0iVwAvo9aL7qFQScSMXngamE8PqOuk58TwQBVC6hALaOi4F6thTieercNlujgX3zPuX8ewYBaPrQAEA9EHMgqjHHw8F8vOU/ZRa9rIsYTNYh8MQzmHqiYdODj6fDHf5dTRHG9C0G71P9WfkEcDwaGGADotAo8WjEetBHbX8xtx3HoMweIlwfWujDfvvubjhiT8Di1IYr89HCTHjAXhrwWD0rpeRmVay2MxxsiCWGEZzY8UgQnrGcEijHkUwIoGnMlI2QA/Lnx0GF+adFk5HkixoM/FxNVlyIbnc58PrFejBoRoyNL6u/HfOz3BBEDKjGOJ2rRIIciXEKHt/gOYxaNKYKfPZlaGAYGghsOII4nv2tMeuqwM05G7XF0+jNjH5gyUtBajuMJjEE4HAOl1Gkczw3/q/j8TB8wHp8wjifyfJdTxXZEVTy82qMxDuTgGhL9LP2cPxuCtmPvO4+QUMPgQYARqdZiTCGW6ZSE+54XIiAkMtrBtc2AaxwxhEjllGuh1gvz8Q2gdA3TkXtiBJE5P+9ERCDmG3xCle4JXUHPfvCzro+2k51CyT0VUQ+dAu0zK/fPMs25eRU5EaUt9Pm0vRgTGIN/LqfWDjeCyMYIDQoAXhMhaeSFGHw3O3S9EAKB8fhGf5QYxye9J/d0HG/I850ZQu/J3PsHIvJGQ2MC8YYYE0flFXm+f+W16/rQgyUQ2ZAr19mRcOe/ARS9FL37UKRM4Dr54jrwfP6kkV0vek5HjUguVBJm20DJI5zypODBK0H848kNUbriiFzrUmKcTC1Chm7IlUsb5agYDRFtIL2ZlYo+AEobe139O/052ClAKKpG8XO4odfNuJKfcUygmGpU5/3ZB5pIQ9uyFkxH2JEGfEi5N4xXJae7GEEz9fMH6lpEG+YZUk76OmWUgXq905gLWvegA7nOdiZ5vTOVcCqgVENRQa94EYUAyNe3/Kv5ABajWa2FWl8Y4ZOotdZJpKO0oJS+Aq8OYMCgA7SdCkrj+ujvQyXfu5bg9UPBhGipzneM+SD6CqagkQt1vqNq8d2qkPmOYrhQ+jKBdSK17wxiEzHtIBTtc+n7uQ44i+g1AlUXkU5mp+bIpSAr5yHbLQWAPN911l6Ie3pmDkXvXbbJUkpkBJzJ1Ez2SCesVC2mbFEOySjDTspIaK04ZhzKi06MKbjzjH0AYiDwAFAYMRV9L3EBXFSYNFPUdnRJYBv1mAAGhiLxGKu9XkctRazA4CbFBEb1S5i4wnj0gff/2njDmwuv/lAaI8MXF0OuYzUURDDXLZQWeuoN5G+zgMjO7bU7GxXLeMfjkw6rDHYOGcNoZ8INKG3a0jsUCctaRAnP7/C7KgnPjwcNfV1tlEx/GI12mqbXxo56dmSVF6IEVzuXH71G9LUiO8PGS+cyHp8234DaEDrIBUR/cWgfA2g+63P/uwMMt9qR7QEvJLmdo5Gi0WGul1DJtjE8PqPWiXl8QmrPo8g3xFBQ8oEj6QfUwnw8+MyZ5MbGo4NWrte24eN5Q7UPvcPAPD4jrxcg3ijsJGRvDBhaYSGHjt7inGzrDqzlAKCfEwVLXmRMojOnunL+DIYLNZzOCglc4ojseCJQN1sr2dkwL1GJ4TNjNNFUggjPMWq04UPRQIcPzrsBwtLhvCY7z6xcqBIhJBa2HBldAQmS9GbhyxAXIJJQJDF8tpdsQhPoKA8oj67VsMkcCwx/i88BMF80cx4AkY9yNeLg0VHMKAG1o3w5QthpDkJmGseCF8ibEMdTkC+AQTJpmACt5WpL/72fazhdkqGM403oIrczWJds0amcYOr1AqB/T753XS+hQe8NdhSrGylXBRNvBDNap/TvovP87aAuY6jeKx7KbMdPh0dOx3sRcew0oG5OuJJppH4OEdsm1ouf52dpzue+Z7WRouxjv/ctrTC/oAPQz2Ci9xbl9xnQM6KAKO6pUqMdcnOvo+1V6RV+1Vkg76fv7M/dqXoZVd3sOJp38PPajk7tiz7Pa6LA57NoO+50UfY45NBLZ7sccHw2ZR9jvimFHjhQKYMDvVcueSu/tz3MhsfA5jVI/DCvHOOxEYCiOH9uCIA4YpAkM0E0xhtiPJAdNU/E8cZqA04scNECDx68dQHBfDOOsTkDEJLHfGjT+cxD3IeJHNycBQ2ELLwJLPMcY7519C6RuchSxcDRIfi8Th2EelgReMeumJlTyJ0e2EjMko8HYsqrN2ehffHnmFyuUBSXA5gPjDH4vJPvN9++i3x9IdyWkZKJH4hMst4IjPlkpOwDdvQ6QAiP5OmTP2vn6OpJ6r2NBmOI0KSBViOVUNTi4RnzQGZijAfS6dgSAgRu6MV7LsRp1ASIEyimijqoropxrSYRZAxE1g4U5d89FI2XoPfsVJUIVbYe1RHafz/i6GhMBOS8X85rCBmNAzVPAKBN2wG3bzkEzr3nJLf9mVW0/3G8ia8yt2cCW5yQ3oeBhfY45nO/V5B8bmQi5DNUQAgEMhPz8SAvqIBVeSFy4chKxLqY99WHjPfSAoiM4R+yFj1jRwFgIwl5p7zeueljNFtfiibLh+j1zgeWoWW+gHXSqK+Pzg2Xy37rhAqd2xvn6ghTInYYoRZiXsjzQ8RlYX38CioX8nphvn23vXMcb+JFTuB6Fyqmca6PH9y88tmLBhRiTUH6G+K5Xjy8OoAu76aiBBBYqYqQSqViRTrK5frS68Vy2o4stXKnJXkhj2yDYGR4KScm0hrzgevbv7Hz1gg5BPC9zMMASPEclRdJQ31urlPvJD5jXVh6r34uR2JHT61BR0WA75oXS9hgSTevdyRY2l0vpZSq5pgILzuw5rZ2JCcxLMcSsfdGwarRwTqZBgEomCc4FElPRCqqFgMj7eSDNtxrtglsFC2x1qV3etMiXrRjgGXKtYAxUOuFPN+R5xft40Y92zlUl95Z7lw6by80/4RgxXHxO+bzG6zziwLAIY5j8RytF1HuOnF9+Zu3PUiMQ4gtNlJd10uVsEBd71guf8vuxSuFcTrt5hbNOiKsXbKskyRSrVPvSsMqgMjgemGa9xCEdwSqSkQN6Sr09wUuEkoRi7xJ6e8aYpmYXK9eZD5b9jNgTBGLJ7D0e+U3C+WD0iiko5KRTLWBQ7yA68wQ6VlZRFmViMdz8yfK+cIaB5dUZQT8Xf190vAJI314oMPGZy4IOq47DyG9SyOo0WiFpV2lBCZIsaNHp4ZCdia3AtVIzrqBtoFOPdCIaR++1VULVlReQh4nupQ6qgk6vWATrVz2Dzp1Hc7N3VxAvqHWO/99TASAxOrobcOvuDZ8vjYa6edvG64OVu38r1cjsjRJKkdXuYAlvUQMYMle5+Y1WLm5vl4X/53tQcgqTSZL98A9y9a7lIlQcVUWf9W6RJC7OjKIxErnSiR+QWd0TKDINRZ4rujIFNwLnaZ3haZLtyz9cv/keJxsCgFVJo6oUSOkUGsVJH9omElWfhiPz4RGEqiEmNqhnGY+PjMXsoEdF+bzG61lthd2pAmRKS5ZjXgQLt55i4NOiLXxQoy4LTz/vdOQyiZpoysALyCUkmSyBCbCjJ+DRip0YPyOjYgEp2++q9aFOl9gTVqltLWYQqydnpRIUawL8Xhro4gYiDJMfCDz2gdNhkdOQuRiV1HQTHzYEfUxUcpX5WRC+fJUypN0VpBTGAe5YwuJXHlRdaVTTzsYk5HHE7UGUyoASO3DEGgXTM+R7eCqgJomuRnNcCT5HKi0OQ7kGtIlaO1jp2TxEGKoamKdqdvBAHO9iOocmLQm45gkPJWfVwHx2CXncbwBY9KOxwMxiypfr6xQyTg+A3nKub6hQshZu4FQZK5E5cToqlsQwcphMV0qjHgoyEzEPJCXkFPS/sbxJlLWnAbT15Jew+V860LaUYI0QhxPksHHg8jRQd8BDxN16vkP2or5K0QgihxdruygeUSMYDlpwzV7zDieXDMfvLz2AU1CHsMz5leCua7fq37OA5w7CmqDYz4FUCzYYuUESjVC3jxcBooH/E8VpC6F6s4SN+XFkiqwmfH5wJiB9fq2BUZU5IFREdrUcL05fNxoBMeu3yNUrZAKMAb1E7FsGK4GxXZ4cwuYyIeMrYw1elAUNp/TP+sDx1NG/gUgigo0ow2oQgGg8ux0in/+aIFZWPMgJ+IDvJ2GncQD8/FZ5UqTqe88uM2hZD9TSV3K9PLZ6U/EZCoWofyZVYmO3Nj6GD/bFqxFr1sKVYa0IltfEJ0y5/nO1DOm7IopwzCPFIPlVacUJiszO2ChhF7080NlV1gvUim7T8zHZ1SRc6E69EU7HIrWmbCWxgh0PD71upGbMN9xyeeolD1s8+KNrOIt6yIoshuH3qXDWdzK2tXrar4sYlI5CzCQSYQ35hsSH51G+h8HzQjqLGrAnIO939lESXskqe4iFiOUGWZF3spFnqBUjquFdb7jePsuIZ5ltipZ8r9vysxQijJdPhV8SnrUeLwperjkZOJxw8EuMWW2MaBI7jQ87xJawNWXJuUkiBo29hFAEq4xj2W6ZDnzON62UWiBvypHzQcPSNDJjsenW3oRnYaQzNJrrdc+oNNlzoF50Gitp6DeRGjiJrriWpRg/Tb8MQ44+4JSKsuwTfaTeLvzAUqhbBt8wDb2UuqS1pKIaN2pxYUq8l/kb2jMub5teE0EUY1e6zo7nSqnFBKu2WlafFbiVHCM7fiK1aO8Vcxal2EEacVquYUlZaNn94u4bG+ex86vKhGHZPavL4j5QJb2pABXFP28PE/Zoq/C1dDfQbEUaJwieA3RDtSOBaAu5oV4mkEYTWJCpH3mS/5Djrzxj3iSYiB2cHF5esw3kaEiZVOO/RhAPOqoypEXPQpl5DJIkU3DhjJ5MAvAen27kUOuJup88JsUsnErNyPcerXxVV4ica6OOhDZZg7AB7N7F9L6irMJxpJYzDkno8yXvbkY/V5DRlN5bYitqkyqGpLY4m0bJL9j6zVKuWOX03S4Etgl43Uiq5oIWx/fb0dX1wsZX/qQsxLDyLJe36q56S5Gqr0OAIYOKJvT1naQJs3yAuohopVIo9ZrH9KLaGSdXxQ9r/68NEk6DvFJIoKTVap8fcE4tmDrXopU01anS0BRVNROlIcoz3cMhFh3VS9yYXwVERkx7cTNy6zXF7jxCQWS0RIGYmweIZM9OUTIgugRQF3I8wX3eVQf2ot6o+PBvP/kO8OcTO+riE+XgiHVbebe9xDpvYRORIi2lmisXrfx+IZOyk5Je5jrwpjel6Mb3ioXcAnlVGGpl6rWhQId3JiWmX/IeX3AFZbKk/0mogwCHy30qnWh4tVEKs/XC5FnHCNGIXaJJ2oC0xp7wZp5NIwEsMVYMZhfzSc9oMpNzhFxACMm4vjcEX0+v7O5AEBlzUc30KAKFZsURQzM53fJVTR0BZBPjCfFMSXugM4lMJ7fMP8UI8xIBHSt39BqMu3I8wvG43MbLfNINm7FpFGWvnsMQrwU5OwcWVFsjAcw34BK8ZkPDITk8jfJMfZ6um9lPCjfnSHhWjy4hoKVYyQwn4p80UIjVq0AC57y+kAcU8glen3zJJnZFYHFahWrEy+MX6Vwrbwwlb/XOFCLKV08Rx/CXYaDEId4iXApU2KiovjKAj/b3LAzcoXKhHO3BzCVwHp1qrTTLXaiUiFcYGPpQSenFBS3d9oksCsyUFpzfG3XTs2mOZaHqjR8xzjeMMcDeX7Rmis1m/yuPL9wnbuKMzGOAeBtp31QqTOA+fwOFpxaaR3HgeN4wzg+KeAydY7B6l3IDuykgQFMYM4nUhJ2gKXarBdifup3j/mmo/TYgRZKrcfBcyKkzO8CMI46NsNOZNBwyaUq1/RpMvSSUPcd1EW5LhTIurvnICuFItQ/khZ/nA2V+a67orE+vi/1HDekCaP1AqDoEOABXy/gVRt+yTDLFZZKdojWUn/HaEjYxNkCEjuN6c9ymdQMfQy45GnSie3ugaxdIoSgsRcfyrdJ+7zQ1QmVzzp1gkqVKq+hdSA0glQ6hqD+g3LrT82LeF3yerWhQQIpdlFKIu33qgRSEQpJZ2t5drlIrYguAvmrzlKRi3WKw3BrQCUQQjsqr9b6EFu/0VfzI66mrUtlutqOByA892HQ+xP33QVWiTFilzEzkUqlXZp3iwFT61RJXV+ShRqy2VBZmB4CFkllfmB2KlaUhqts2yI7IYkKopZhMnuyyS8t9xb66H1DYX18X+kl0I1wev+sD7iJc4sKVQExnxGj+RKL2IgUVtsEEfLYe5WuxEh7Qs8ihOR+FDkusC/poLAdTRJtwsz7aoRRrU1wo5BVYZ2D1QdGTFSo3g3Ceqv2uqpiaWo65700x0BEnfNDPVdnW+oU5C+5RHlLWyLUy3FKtqvIh2DNvGXlKhNJvJXXO2Yw17XD6zxwDPYMoDBSJSZtToWqCICET3KquevkqEJeX9TOLgmyFJkDYH7dQiRCZXf88rNEEKsGXs2CW2glIU6jm0K+ftDEFNedhzyvDzYZ1QIG9zkAfq7RBrCNR6nPGIc6cp2Dn+KlonkoqylpM66ISSOQiymj+1IwKI13lWDc9teaDXeLrtfmLuxohiJqbK6Cz/ixRWduhnJ52KVtlfxboh1TqZmewWI9UO7N4Fk8QHIOdLrqNcmLqZgdYVdi5Moz6eD0cz5rjvLkYRbCwSOeKKFDl9c79bXd1Q5EdoIsAV+NFvr5YqPEqsSoRwdFpzckd+VorhficD1MQS4C6/VtHFhncK7BAsBOzq3mA5nT4BAQuFfetepftUh1faCOTxuVmEV2peL82ORZLiBWQ6/26MqXofkUEFyWH+ko3u2+YHefjZfVlomh8lWWG2cuVTC4gd3SHVb85W2jjSSO3gxYqotdajSLT7KfVYxxS5+GSlxjPBtBsKZNRDNUqXFJlQhhIqYrTux7qFxCdGg00KhClYn+bzv4XEBwy4ccg7tsy05Gzp9ksA56S7K5fz50SIh8VVqydmOW4XA3IV2vjmQ+hPfv8+yOr4hAITETvFVJpCWUxWj52NxMAZZp12s051M42xHYWUc99lwHR10UBUxD6G9xtkddL7QOAnaCEBciRHh+8N0v6354NoxYqxbndKwLMUjIZo6v3nOMh4hIkuzZeiQ7gVBKRQ4JgDg6BUU7O/FATHOzPz+G0zlpVcI24yqdqmE9fqHgqqMdiLvN1S8iUXcxf/EG3mWqUdi5JFheRHtrl0yHqgSPNs5wxHVvRfEBLUUNyWz9YP7ZGIfgpEpK44FN4+8Dsdl5QfbSiyD087GfV9/TUUYtyt0ibQc0n/v3usKgv5Nz4AF/7hLsfGqhp/QQcjZ2LC5VYngKlDQtHAST5/t+/k4JQQ2CDt9OVRy1j434bsbFdac+I8aDqYrLgzGJKmBNhfgLf76rC1m9p47S3sOIow/3OJ7bRloi7fU9+hB0M9h4bGjvtFCOLVobSIl9QOVl/RmKXNBQo1WvlVoM2nnIJo06ms9xancjTTv43J93PLo9e7+bnjl3R2b/PlRmDDeaZTtN83iO2hQ7SWMTErThJurq5A87PZW2JmQPDFrokrRL2LvFnBLwIdu891rdz4O5O6f6vYey8RDtMIRYfQ6OPiwBAK5zb+04IjCPb7aMOy+4A4/OpHZ+jp3PegPHOJS2EAISUsuJhJRtjuddAvIshBOufxvBcO7F2ghEaUpFNvFlmNjVhN4codDiXAWXMBuCOzUSudnR0S3ktT8jzy8kEONSDniJhdahcAnN3IByaRgOy/ubqGxHPcXKO/ICXS5ueXsmbjOGYB2AoWOnh+1Uq1FhaGJWdzrCefTYlQiXC60aFcNf60Q8PvfztxHqXQrYuoQwx1FtE2M+u9muUkaOjaJYWrxpVOZBNDKo1WgUN+jw0pLydnjY7938h/UKNPiSrN8lZx7sB6s35bpeOJpuZ0p4tB3ILV1GbOKdaPPaAbYRiJ7J76D/BkoVDqHase29qmTDEgvCzzA3J4PqKiID+6vtugPA3Q6cxiTgSWmEP5sct40ah6g3pFcRJjEjjj70/G8RU7248lQ3LqMj2+Eoe9vsYI045lNRINoZtNf2IjefUXwez5SIuP384uc1SVaCZVP7ub56rvuUJebtr19z+O1g/H29eSIKOwzBB8cybKnqTCr5+5QLsm5/dV5tY7fWglHaRN2lvzu/et64OyvoMQAYHez8dbYjpOPR+zR5veXOnf8XuHbKyduBKCrf+aIdae9p2Ghkw7Rk7nVzWskIsdHHOmlfQfTg9zIy3RzZRkA2/OEIKLRmlWTbpXmAjrpeSjdfeSLZTfDUvNOOuj74qLx9p9r4x8Fy+TgavXS0x37WcFpwIxCZBsuZSWfEQVIaKqRU1ut+R40lohF9BqDu4m2a/h4GqewgwJTS5W07kdWIkfa4u7WNwqA0k2dm4UCMYl/GpRKWmGaXneJgTqRaMI3G8prR81icZ+6ORZdU+bJ5fWA+voH78AuUzXrs3l4YaMMBqzK38VQTlxtKi9DB2gsX9zRksHb++MTKhY1EGolemPFARClajT7YPlR7pkDdDvKxyTmRlBTB8OfH5IQr8xs+zC5R9fQxHUZ3B9K+gxJyyfCpFdFhnvfWe7dNy5m4YnFLpzg7kzMdWNrl4VrrBGq3IjuN4D4qgOTi3IYwNhvbALHhTetCdMh6Toj6dZwO+FDrePSfpSsNMRGS+JuoRAweQ/EI++AU5nyDJ2UFqoVsvyZ1Dga+bv/X0Yb5FqUesIOLADuhT5bPMeDmuFaaVgHzwIhjk9R9Bogm43jofHq9sAPY7Xvd3v9r/nElypPELM6COmJvP8cU6Angha/GNdyqcnx27wvPutXMqEDUsYNFSBhIArgOrDPyfKfW/XwHUO2ZuOnkIfLFKUJYrFosDXqxF8wq5OtbMtiKrhyW8mzPXuNSykJFm50Cyc2dzzpKu4ybyRFyrHoQurbiL400HOUOWL6Lu0dPToVqmAqRO0MbArLNY76BA2FcI99S5nDECBNHMqgeKKxtdD1b0XiXxbTwQgKMrjvyz8dnQu6L0bdzT3Mprq8bzZWhuduVB9zp2Hl8R8zZ0ZCOMhAVt88pEalMx+pS6bOjUnUaSmevKVRjItdHP0skA4UJyQ/ajIYAACAASURBVD3jgm0JfKghp3+o2UqpVbLhCSLYOzXQ4dvCqN0zUjo+LkmPUoUlAhwKn9sZX7mDYQwJkyYwn6jrxHKzmzRGgQtLP0OSN1XRkEBxqSypvpomQHPbNytwQnRxt9PZPwucvYfh2ZqD6QzPyNj/n0up/Eb/fp+QLYwbQvMovt2xvBDx2MEYtp24na8bunMgiYmjqqJ17wF4DkNPUKpqlV1DE3XdhcnLiBtLXQrsow8hF8mHcqMIpYEwixv++YZ1+vji33mx2B7OaJvrnfB36MAbGZjVDuy8LJe8sXgVeeO0cMslz5KepKy94LOWuxz1DOP4xJb6W1m2YqcjLoGy3PWGrHdFBCDPbzEVXTwJe0npmNc7hoRdhcLQuneH5DoxHjdyLGe/T3M9mj7VytL1RTnqbWwAoL1+dOrYvI2JQqdr+p0BNMdDB7Z1Bt7fUOrp6oshcn/mba97/KDRpaNkaxGwOz/DfQqbB+lmQfFC5mGYijHvH8cbPyOIPhrqKyiO8RRTcnsepZwBAlX283jeKrt43Zlp/iGMeABEkX8xB7Znk2I7hLo5/dtwI/ddRRWqXu0MPJekhIpb1SqbJZLMW/AqxJLKWqMQeb5fcIUzPAv2xrPl3D1E7sSO9RpHCJ7RR7l9O+GJwp6M5JwnwJzeughD16GUgiSNh5OOHZ0aNEXn2R7Vb31HdrnnYEQw+Wk1qYlTHjegcqvu7GEVBWL2HRRwtSNzIQbRgLUZmWT2x3wCU5Gg1G1Zg1GniS9+xjw+weP9nSaMTlEgGPfY8x/12+NgVIIERC53zcceTdcdhY4ctfY7KYcc47Mi4lsb9Ta2iVw7B7bIzSlBV35otYh47IPfbL6Ms5ZSJr7bUJnXiMnBo9uqcRPz3Dmj5jm2I2iNgj1CoLUl3Q6gUXqeUQH1ori9HEIxdiz88yWnov4b63eqgGK7wrjxCCS2r9Za4P55jthWgd5UpMx2q59na2MCdS0G29xiPadfLghYoFUllezxlJOWA9IoQAeNnjeRCxXZttPkfQqNWsyoYNCDt53OjikwnZjqhMbYVatyZ63TMK0DxqMOxKz7nMDKpenJyuWUe3ImAiW7PqBdKnVDynyyDt+XvHCh5vGJTsFdpGMCS1FC92EQPj3ZP6IIaynuOr+Fa/38/ack4VOHyRBqYC1O9faoOqZCn9CNbMVy1NDGzjiEnMSuI8RfHFB3FY1PQpah9+8p4UYtoPae8ybVBOVnnG+SzBudTSz3dgTbv8M1cuwUhajKebeMWptrkrc7XJvQo+PKPDHnN4yu1wdMzlnSPo5PWOcPaIza6+7Rcd7tNv7uBLZOxHm5yeMS7yGniyA0r2pn2USsUyHxQIkX5uMz1vnOINWlvQHo3hOSrQFPE5ua3ZpwhWwqx7kRl0oRnUoXXrdnJ/M/FGDGeEMO3bMiBS4Qey/syCWO60hs3gLR6zHmgRpXI55QUPBgnEZCMTAOytKrgBEHoP+m82e60BoMp6OaiQKgCwZRhVI7RKelWofuuRoKd8Wfm8dn9HUHeRtTGe5SfWP6P9/ktGcdqIqeFCxmt2BxEtDDU1Sa6k7QLs8kstSIsk5eflJtQgDQarQWsRjejO31uxvTKEGMPqPVhIeMBm7lnUDnnQ3f5AzYNOaGr9Uphom2lEDM8LmWqyPR6QnkgbtkLA4hLQBSZGllabfhGyZrvsQ6pfa8dRcaZtPUaBDTRNfVzpLVBQ1x0YHL6wPz+R0K5QCRu67AXP2sdX208ZREdanDtc4v4JSy95594OpEl6Ydjcv8wwLqQ58rp3Vj2HNJdTg4yMglSJaxP3C8fY/pmWaEQmrCjFcj2Iqz1z3MMYf+Ww1d68UGvO4N6aoDy51NX/rP0pFWTi+lohWy8RRxz0htYtsS9zHx1WyJWdp/VxTQdpuaEVGebJ+LKUJZYuDUMdUqwACWbhA83nqfgYW8pE7uNOsSUem5ria0Ac/ThJxziB5oG3ayFU5Fhi6LMv/h8r16pEAZPfcxybCN2DC3hRyFrxSOJhV7AvG8CVhUqybiINs/5qMbejbB5jseLMzxS+duJLtBP0PCr0QqgsN86Zt4ymSmbntyeazVmXZ+PqCuGBj2+28VYe9lUENqO5BQKmHU0TqS9uyUOX9V+nWZ0PqUJrOEJgxlw+VJ7J/XevjCGioy0bl5l/xwLzFvdt5/3kORhwRkKjn7Pfa6KFrKsMZ87jLq8B0oTBF7XkMMjNi6BdsUlFLNg2g1jOpidvrXIqj5RAuGlMK1wGls9GsEM443jPnWDXNDiPCr1MTcicq+dtStsTg+bTSj/4ajshrwADVEOpUwHyQ0a4KwD7vs5Y5yerIad6VTAv7B/n3vwU7JSLYzft10SeYrjGw7/UMHu8AmwCGCGkKWXcq/O0ftumeF9PiHWgCqDnsoTui13n6TRySFNoN8PzAdhRTtSxGvv6yqjaZ1BEh1wulKNgARLnuKKwkbuL9pM8jkQXb/ise2byFSfLVwLi0SQSgfLPDaQTBi5VqYx2G/oIXyM22ibaceEENfOlcizjyBOX/VtPIWKLkun9sBOt2LiRjO/13DF1Hb6OZWcotQ+i/jCRO3pYPDQ5Um2cChKMy3C5twhA4K4KlIdkiVJxHC1GEu/jyVlDowbfyFGlOT0twKLVSIyy5WCEsg363nSSk4l1JQu8zSK2j5uTMRQTstkZZ8B1ccUvfZ7pmWthemd+YvdgDowT3r1EHfE9mhNC8U+KAxi3QmCobjAPKGiCDVcIncB75u0otD0duduSofr1efJ2tZYNvvigxkZ/x7O6tcH31WCiZ4yZ0ETzDcxxP+fAcGp5XhAsGxbTQGPBT4qLXEum4OwFCpa7Rj0oEsXxRk5l2GMqZuV7U0OHl58roQs1r952lNvu80sSdKwyKlZOPTOD7BMu9cHzKihaohKM5BOD0ApQAMz4Wg0ae6It0cdG/Qai1/pW6yMvTWAuUtFXP0F3HmEmg8vmlizOW6UVIyjolcq2eM9gVIuXSuNUdR5FI6ZdDa+J7Se/4MP2Net7suy60sfJZhcVpivb6vn2HjWK2P7eTG3INmUD1blenkCzntZICvFJ9dpVDUAghVPa8iEvX6VhGNzX68XpIpqkfe7ZQx22h3F66+MzjvZI+oY3TkFYqKilOlYgA9g0Nsf6fNs3oNdzfq6giLQCPRjhhVqHxJqfum96d9Ik9VlpwWvqMJ3GSPlPcqxmxqvzU8ij7uREaSODXH4fGBClu7KdKpzjoZlD3/pasiTrturRB2mHLOYx6sgrQ0IG7B3AiEymGrcSsvYC0cwxcQ31hskdOEis5VO8IL2oVLX9xYxJBz4Pj8vvjlrrDzhvDokdSB5K7qVOWtVWR2nSuPon7CJA4j4UUxjGcKOsURW09txmf4Mt/SodosssedMYcecWDVuaG97q9sJCVNQsPSwaYmro9KtCIg92wPlaV0IO6Hwd49xh7H33ltCMYeb1jnFyGSJyJWO/UxfHGOIgxunJMi39QcR6/78J2ZnjE6XRUSGRxEL+zDeCJxdjrDCPM1CThCIwe+Ij1JxOX1DispCejcDpCNPCIGm7madH6q7L7tpG1OhLkntlsTAEQP7xlh+fgehUB0d7Rdc6Pu6Zsv9AH3sSQjGIHAxDw+wxDezwYjxE7N9qGKoZYGlbDNk3DPZFdLjV+Lz1yDcvfuJykgjqNL6nNyKjovLn/xc2JXtkqonN2rJswZoNgecQkRctzEGM9GuSVyn4s8uqTc1x5CZ47zLNARVrR1R4wRey4BIzNgWXapm7SHjsaBym/376c8vQ6BYREA3DmCXmSjmiXSVBOehlKcMUuLb0hXwJCWIXi3QusfIFLVhCDe5a05G8OluJhPdjYq0lW3KocEagmLlRitXVqayPNbMsaV4P0ggraPG9eh/8/1gofOmJ3OpVvGL18diZ23dsTlc6WM1VAT2FOz2Gq/Ou1h1qFIaxm6+mAahclQckmRWxr7rjSngiI7E9T8vpciswRVCBT4+ePxmZFW6YAd1J75ICm5uCkUUaoVtDsxiTbYQmLgsdMxIYuuMMTAOr/lUOmxmwQhXqIZ/kxouMRXPSAUy71QFw9GZjIDtENL74UDxi5Bx41shlCo9QhMv91zw0u4xnhoQrk0OqX/TxPOAz1lS4UA3ka2L3uKwQlquT6atHT66fVF6fY1jRWwDIA28d7OkefOIw3jNn1uT+Xyexj1Y73GkeusOL/QG9dJ+K+8l5DGpB8fMPG6HXAz0WLXdejoOF5iXA+l5Qsx1ONgljjdC+IzUvLsN72Fy4vO99RRuXv2nRqoxOX/7oXJ5iu+Jm8WIu7EqR3h1boCRqCl0pcGyYSmHnXKdZvx2fLxezchesFJcmpAUCivNUTNCwHlynJIfB8ak8u7TDdu6+gc+mbgRopujjMRd3cosILVzjAG0vNK7cjXuZGEIo95k55sNWYPGwL2LJBlAVm5D8cwnn0Imby3s4faKKLBuXltZ1e3Pa682BHOR6RjikGlJTyiQGjZFS2l00vPYZ7Ie9S3o9cd8rNMmy7b351BK0k5Y6R5LKd0qrwYgXtPEqD8wCg9qvfCh95TuTyR3c7VnEm3WDgohz89KNTKrW/pQoWQNFTqZVPf7KBpfrK7nEMT69ZOOysXjjFmUL05u/HrXmFgHV5lv87XpY+I0aP1Y3Ax0A4ELTvltGY0cuneBr9o6FYkzchAbVmuo83Q0Nz74YbIJwzr2amVON6+i+vj+9ygKnZTNq3hGRV8VhrY6gnQJFehTSlEaHiuoadJQexJ2+RKpBaMA65VQ5uUkf3cTJGY5+0b3LJ7Jfi9qkDFrkANcF7lwEAN35Z29g1ZgVsJrkrLdvCONk3mapkwsg8yGwddLi6pFJWONCqUw2tZvQfBbuLZqSp/BxTpxZ7tUXcnFkBgSjkpGKwyJezU4KqDbGQaTT6+sk9XlvrmrWmpc30VvPjV0suMXRpk6vtEJdO9cWsJ6BYBHW52U8sm9bsYdPzh4gCACFYEXeIvTbPyeUjLDuzepEaG2vApxnpSEJgLFZLiq9UA+qy+DhHS2yi1zlugirZx7L0Pjx44ey2t92FKsBDzM20yQv/9qLFLn+6/V57ocpPVcmUi0tr8uEXvDW1dNu1/hkpkx1tPwxZe7byV5aGganLceugFa3eJ8N7xCexeB3XZCb5zoLCZaGsVjjYilya7vOqSbZOJo383bJSCuB2xHKGMgr4ix/z4G7FAh97HrtGbo53W03LlnvzllMvOyp+HLRV2BG2nNjSbwA7Ia73N5vZPtZH7oJv9b9QxNI/B/I333AbYTl3lQEcjo4leyV7RW8/QrcNSTYYsrTpVva2BS6wdHNTcZ4c55u6LaAeHbY9+dfUO3fe0Je8qjbZtaX08DdulVo5eQAc68ypf9eA4NRVf12eosPkAl5hN3sqG8vpo1BSOdL2P6ANuZ91q5Rb0bYdWtskC7PDv+pCvSrptSzc7UXA+1vkecX5R96fYbeXYWC8sQTR7Y4AlrLw+MOpNfMKbovrHhn61RHLJcHo0+sLSQlVMRADrJNdBQudsj1dVbFBb77dJQPxsVPVFLxtGqTlo8nq8ofLdwHd4pZyFQnKAMfnOZKU1uVu5o5WMeyTd1ui7OSzCWv3V75k3DiKvd1TwNnYq4b7IZsi/5LkPOS+YFrJA9vicnozdApst4zWCSztzaz0k2TXH0fMZPalaCk5PeI4gj5N566rUnrkeX0of5oMDZCN9iXZtx1LZ1x96HBucQq4Lo2pPLhMp7b6FnlcyH8hT11sO25vezwLBGG2D8/iEEuraKaBGyCkIeKp6NSpwGvUC1MBY+QKSI+yWBVgx+hKt1DsgokfdtWBLFZE62QyY5xdOQV+vJjK7Sc7B1+rbQYeX6wO1Lkx3UVcJyc/bO6N/zhUaRGBUwlO/S5zFnXDOPPcc1EzGUSmXO830PqmUzaFMTHPz+gBe38YxxlEu1/TFJaBk1xHGEdl3lUYlW6wF4Xi42DA1bDgoYD6lszioCZWzOY7PWNcXuOPSUMmTeVqUBZYgkUQ+2wjMIYi5Hb5k+ezUYEgHwLs7qKGYtEZsbcmOZo4GFZKe+/tYoMY8PsECmTBrDPThqnx1RCLBNTiZSjm9EdMYs9V6iF0hquRmjeOpOyw9cekBC+ESL6XAQwarZ0AwFTJBdUsHqhJlROP7IMLaky2oq8pm/rs/QIeZoqgnqqjAHePQjVmvnU+7N2E+6ShcVRNJO4QKhhWzdhbrxBwP8Qmly8oPyn6syfDAowil9xSVhdcf0d/DP9vVGR/or5w86GCN9MbxxHp58LJsUmnj7MnqD3EnTMenL+UpNpDZZp0Oh/iFu5Br2676rSZJ/VYXM3L2e3mNIqPTK17P4J4fVQKhP5dwD9NVraNpgxpCHzPEWbwh1hbk+ZqBAL5Kccb8xM9+f+JA1aAWAChI1mv1nxYsdWgtwnJN1rMBgdyTna4XD4NShoLVoCfbe9M/m0Ku/HvDri5FltBJLkWp2c1b1ekQDWcP/SApQ839qd+5EMN3fdTOLTfRj1YxKgWpuvYGOj82y15b++B23r5pRFC0/8lqAo8fIQKqeFv1ePg+i7tIaisyLbzqKo2UfNYJsHpB1Of7WMbklZKc2qWc1wdnXSi4Rd5VK00/H5P6ABHO3YdCFhFl4k5EX8JVKt7AbgKSqEBVGhNu4HTrbsgfHjBL5McJ1H4eXkZEg34oMr60f35fbG1FXdo6df6qCuLnpbtR/8+U/kaTrPrzbKO6YwNW0/a6HkIvW9m78n2jaCGfygtLFUEgpSU6G8ajEjmrvwOLe8905IBvkvO60xGp/6TTNTSCsnShb9RrGzxQ9dH7694v9HCe/Dqdv58HhIKs5pvo+VZedRSiSOw412In5q7jKn+WV0QVcNxuElOE5D0d7Hqr8wsiAgvnV3k27wjhw4SQjC8qIhln7kIvtQox3zDjQN+W1HMYg2TcOhEl9rnzOUW1eWD64CGA40GWHl+nE0YSrOhoIlMBhVvpWN2MczzbaBy5uaCeyuUNlSG1gG1fptz9GrmnKznKdl6fufdPEbfnOyyKndCcR22yVfNH+d+3+QkIdReyQS5iioyVhHocRI4KEiOe2N3Fep+xLxwievHM1YOir45Gb7unQNF4WOLu/bY9pCJ8Bnh73F1ercFL8xNYxkZDeCgFHfNQY10J2XxiEOnSpvZ6Hk7KwQnaQ9skBxATMZ6IUe3EHEDMt4xuTHsqNf3g5/n5A0JWdKI817U5OQWNzHvXKNNUz7XdArQdeNwwZrSc9dLBFwoDlGqq63XdyFs5WfYLaQ9C7efWqihO0jHZWXnbJa4r4EBl9aZWcZFhJdjXTLe71OxFe1EV7df1pV/SdeR1vTf0bkGWSZQo+CYm5JLC7UGjEZzHIofhEg9qAktE0MpObThCv/YG5IVaarOu1CU5Ury117aEWs9Run6gqET0Qa1lruTq27s5+csE570Md7aRsgz3EDrysB8Ni5G01qlIpm+Xv/badvmrbkQoOaXxFRElFGeJPlhSHLoPw3vJiKYyZC5ORxsTtQrL09stRwcH1qSjrw69GwsZTBcAOi4/ny+/Rm01rG1hyiG2kjHdHLg1NF+VdP1dsdEXbu8IEaTjIN/EKpsdtkvkni5fvVZ9ENapQCpORs8ajSD4O5kXA5LSzxkDS88+hgcakb/JxYju6yhY/RLKzS8wOeyfwbCdpSK+Lg1ve91PnXDwkS24vwNGH/tKCXIyDHx23NTsCC1IlsBrOD810mL1xUCAlZCqCyMGjgDKDzqPTzpEa0c/tw3rgFCyvJWKRAF0ECM8lqw6bybJNBFJki+vL913AOehpQEliviZ9ui+Zt4eeMmZRXvOChOzQ0IU8SaeTC3xFSOIme65ZcTYjWN9ebByvZ44FZ4joQijtn17/PvNYLsNvtprW7+PYMv2kFHt6ovyROtDprkMz0l4Mjol+mcspAtHvFspbN+PMgAcGCnor4oSgggQp6ssRztR4JYv34yKUcLVnpJNVjuHe2fq5pxURSh2MjpQmA+KMXaTmpBgcyitx9lBKaRjaLSbyb6VCJG8i5drO81xP5BSnGli0qgDhPljPFBzKx6dNgSM2AK+/Kfgyl/Bg5yYBkDISY7LlZFG1sEu685Ibm3h/kxUc4IBYOou3BY+yoZK6Ma/6xS9Eep1wbqJGIfmd6xdJKjbvlreAAC6zrGlDOVOVYKBo6rCcHj5AlkfnhZkZC8guoxaGzaPKX7hxCGihF6J0WBoCE66Rb1KwXfX9x214Ju2fXdE/46je8G9K1ToOT/2wJTVeWJDqrQMNrGu903kraWI7nIo2tjd00HYOnfaID0GRUfPVuXxl4MNUVLwtSGkLpoZA3APCPYMDjvYRhB9IGaveamt2lzOGFMwV9FAg2d4mTX1FwPkLHJxqlmuj55F4lvRDLJ5/o1iLkXChcBubbYepC/96VRKJG2radfmnzQMFuJkoqJ/F1XtaAHuU0XJqY2NNiRQ2k4wtjnqz52HV3iAsngB7UNgK1v9e7bPvvFtjFv6tKt4hO8uQV6tdO0Lr8yZVSKS4xRiegCPvisgDmrbLvfjU+9FFQfbGJUV/DvW/hy9P92kl8l+HAsT61ZOHzc7LqAqdlqduSfgjW1HDso0Q00iU5A5sFbsur8hnNtSrRADTPz1Hwh10JC1ic6hpYe3Xp/2ziE1/FWzvxMxHiKFdsOLUkuY/XV6EnUjX5qE1M9nocYeM0YWX2TpzcmFoJXbikPOrjc7Bjfb6sqQFNf9H5Jsz+nBLHILVr+NsZestpMNRXAP9+mft/xWpKOdHiR/b42B1gSK+E2mVvZn7LC100WoAtNIJW+OrBgICk4Xqg2J+bMPyE2FaThvoi2dhtwmnht4+ODZnjxNunyQ0UR1M/b6jLTiNao/27Zge4KY/DBh3ktgx7v1MNserkaz5pwqL5GjFO9BMvFWoK7FdEH74CsIOK8kdPGyRjAONw0S1XCtx22vVDaGpsv1I1dvX+83CoDs8P53tvlKNNgabsGHHHvdHJ0GUdnBrJN34Y6nzultWFUw6+u7jovIIitxIDjNsoUZMalj9xc3VAJYfFRnJwEZqg1+6BD6swoI5d3rbNVnD+Wo3S8fgoqMwtzkMRzB7gupCJdXpwueLAQUotxDAFg81WRhE5HRzgCLzoZzO6KNv1vglS97IpXbr8t9K47SuRhxelWgg5VCIiRmqU1xRWmjr7jdA2pGu9a7yqMJqu6s1zcptVFI8xUSFdFJTeXSOrQWEdnpp5rdNLman6ncVgaXble+ScDvaWBPrLYBy7HuNInzJ8NMPnDb+8XvkWEW0DfL2dmE0hDEjcB0JUpDb+4KRDarAfCUM+jgIxBD1QIpY11695p4Chz3X4cP2BUl37taVrZup0Q0qXNgFJ5XpymBUOcto30H1WJH9AhNw9Ia3GdQxBxCdiAJWjp3ue3Ae+NpcLu1PER4520+qJo8lztTlaaviyT6+aUFmh0AiCjjIKy4H4bY3s+qMJAhr1OHbPByIb64u1aDLy4mvJGCtBgjU12gEutwh9VkA8zjM8fnBUd+RUeZ6NxviMUdk2P1EAMWEttgrCFICW562Es80dO9bvm92+DZ/VlI7MhQgHI795CgYad5iALHAe5ZpE+VKNGow6rCrziM8Wyoy2qNZ21qNkJrIwLkoddeC9fPjZAYWm5ci4YWiXwL3clhbUHAeWpoPdV9qq5UIz7jvD2YR8pGQdlRR++vf+9uuOh8n3J058m+NR0I9K1it70mOuFartpT2uzs0QKiks7msc+M18yITPbQU6SSn2O7c3DjVHdqKXzNJfN4IpJQu8G+emD5kbfmAayMrNcPxE05nYl2bOTkTswHx9b5rI2pgBeTLRbALf2A/lxj+EIzOrzaciDQ/g/c0x1KvHmBGAO6hVkycFhJiigMbF0PzFkQddZRWYH1AmxMsSsXfelI7BvBykx+XggcTYv1tGDlrOYgCOfFNl8fsODHeXvm6iYpwtXr1nrNQ8yhJK5zT2S9mAIhWn1G1ln1ehuHT3eGrsDwXRTP9sp83ttIPyEVL3b5WUz2lknYq0nUXF9klLhFeb/jJtMKu0fEfMqeHJadCbqU7OaqPb0sv4b8laioNu4AiHoqb3V5TS+fO2VElbQZnIu6cu8bHZs/x5/hTslESD8ApU51fdC55dpiL0SrQ+2YWbV4k+3sZ/AoRl/7sIKT1v3c3pPO/4WS2kYSKFAhyUZHUCmaF3yXSXMQBbQa1NWHqiYlez6HxgCQe3kh1sDQ7+T1rhL0aEVn6rnohKTOVGcxWoIAcRlH23jfjl4becFpV4xtB7Xk+0bzMbb5ytpCv34n815y3JVKq1wy5ZUPFgcKL3SQgaokJFujuaMjxqwYz44KJKEM62Z/aQxP0fFlQtv70CM+MIbhv/USippxIGOTdm4pt1gk7lwIWLEYN6J0SBk5DIHHA0iqNVk44WH27EdG90CXrcbzBvvNHr9jHG6tNm9RO+UpMe63/Hxr/He6wD/XjefrUhmPh5gcgNIy8THMY1lbN89Dg/HUowloLgGKArYok8jVDo4IRV2lWhdG11tVqhhRmGHyuRlR2T3bTjM4W6TLt7ilHaoKNbNfiu9xwDNFIyYnj3WPyMA4FCkVwWGUgj0vlQf1CZQb4zZpt9l/34UrWC3eax7foNxiHxNjWmLOlNj7M4L3rGa+Ok0o2ZCHPnkt72Qez8LB8rM+k5zJB1q3M0J8ndCQz4pskm0Q5qC2fijGmxDNoYChGaBgMxg8t2Waaxq9HkZQASNdfSZc6h2NNvdUfYnUnBLFwL6BcPQzx3hjK/vdGfa5BI7NL8jzVv2qPFDeHHYeyldxy6uCY+W4RhKZ+JDp99G6ADQxyWi71YHuGqx87eRCUbjOd1iJaH1E4pL35YL1zECp0yxHrjw3+9+XrjjKx7oHVQAAIABJREFUakSdh9/mQkyTclrsGE2ONTkY0is4f61Npu31q45WvF39AjptiEYW/Di3FVe/Cw1axKr7BUQ4epLWVyU4wcYtmZ+bCJSJZZ63QynSuQqrfDfHjj7cM2lR1O247xjZ62zHUvCoQrekC6lg80++B9eK1Vwv8IZyDwa6KRHdru8p1nFX3tJuOPX6YLkwdsu/nbAdXnRqTC4iPVHKxHzt32obN/pribqHVIN224I9NzHyXhrfEdJl/E5btDcAcLuXl59XvU+be/DkMk7n3nsZfa5KE9/cJ0KbONsJ9DmrpSE6nuqmkmgmgHUjj5UyabxhxNHakSPXFSMXCrdFEwzL9bF7PXQ7UqmZaY98IwmTmrHAttxN2JmB5UU+n3qzmSIUPG/xrrkwiVmVvJZgOXeSkXrjYSilhjHX7Ke+30NfcvZnlyOMoPoWiI0+IJ5Q1A4TAXe1liXneSLmJ5G9diCUTJcjsprSGqIrOvL+0wu4zQ/t9dVnkYX/2MSnnXrdVKKC1xZ3NRJKluAMpZGXmva+LntyNBzkANDp07q+9Puj3y62k6ml8LmrGzS8c7cIqFKUl5rCYC5MJXKXBGsh4oGqF9L6gMH0Np0KXZpl4qnTHlMgktRpQOXiWLrlIEAHnNcXPedNaOfUqRI4PrWzb3Fd0GlxLMAt+leJI6nbgSz0vSM6oSF+IJPhwRqgKMguWW30aIQe7MRDg26W7NF5e+AvByG9+izt87gnwpcDlR28y+L63LxM6pP4TFMOsj2mIdvmAgPHGG6B3QIsD8jYFZLReVL/tw5YG5ONGIoN4hoclVHrNvtigo1TBQQfhFFB3z8YxfqKQ2BHdke+okE0KXu8EUoL0VgL/xWplqf6VoiAvIFA7Np5WHKrm8jiBum8IRBsFUKwVqPyAo7PjDBa/IC6Nh2Fu4swxCsMIRsjkGM3YiEaZhOObuTXHAaA6fHx2liSrpQmjxhsJLsx+T3jQ/MqOC/01C3qwPQME+W/Jl4rnSpBKZ70Ayoxjji6W3dXkB6ouHjdJXwV3qn1/VUwe0Q7lc0z+Dt5cMIOU6lgl7j983JMDKhLKbWOYdvxxIhE6Z7a+yHsi5zkLAcI/0dMZFAzhFxc8/QcTrSd0Y6JRkxUQmjC0/ONeNhOcMrmdgNk2xM8F7dPlRDGBax9N3FEQIP693mx/F7kZ9zRjRAfVyW7gpWNtCcRbi4+gxDRkbkw8gJGy3P0hY545iQm7s1FDcEATbyScg3jK2EJik1E6/oAc/t9/2N3X3Yd/5LAxLJvjsGjfYhgO7ZWwNGE1rCQkbvZrLbgyWXL1ndMX+nmIblbyOI2Xa7Bsq+FuzkLFxAH25Afn9vISjVvNzjFsGDG05feSJxJGswtzEZEFsJxnOBLkU0NVZ3OUXqLdWI+PsPTqPP8gAlfQ+YWO93fCdk9Eyw/0xmsU92Q60LgBIPfseXK60TEJdvgIbRUm8yxBs4icK0f0GiVpqX3Ni/kFUBYDHZ3wikHm1ua3chDpG5Zxp9KnRR9M9A3dZXuEbnpKHJ9IModv4/9nSo9V1G+7TEFnmx/R3hsbqMNZC4cj296Mhxu8B8x1Ea/qJp0IHJ60KP/1D/jQb9NSnJl+q6eiLYnBN87NZUsfCetv/eGJokc1Eahz+gWAgse8z7qUGcxZe+e7qXzw5R9xTHnW0bfSsUPd9s5XC1AbUcCGm2TNxqDFwiM+bkRQMvEQ+P7Y7Z3M7S/Tw6icEhRGDvSwJWJoHdH8XqBhKOLdAE68I6KJrs6R+zoMzsSQn2QzdNUckzaeNPhQ6/D8Gh4b+ktKloH4Yhe5Z4THvip9XXp14pDxKOrId0ZqHKff5aIQ8RX3KKgolnIWE3c8k3NLRytJ5iT91lYcLWf18NqdkQn71BCT/uC5sqTQi2TY2CkTDntoXs+HGxCNpLYZHYjEfFWllND0n4jqcyT8ux1Sa7vy6UfO5+XjY3jEyKPltBbUr4l1+oRcnu4HNmY4kZiYkT1786xkVqEKw8P4Nas1T0XLZdWY9d8skdK9mEpfqcmRqulJrDaitmet6nyac9ptf1qT1BbTg6fA5PvzVVpapjTr1CJ2jbhmS5KjzmXg3jGcu9cG4VXRB0+/Bi7ouAoGio9NcRDoO8ncN6ord4DaaIhr8IhkNIk5JKz8G+RhKy8kDM3atHL9Lj/XFsc0/mglHmO/CLI1vUFlmTTE78jHp87F8U9j54hxLOHvWQTiWgj80HK232SREOE0h1lab7YiwJYDzDmA8t5qdag8kTkbINuZWBegqAqwVVJ2FTawMDxGN2FaoduzM3cuMBBQny2BHaJ2tzJ0gW6EfuQzz3zwRPRtwTd6IZ8BRvSbpcJOZWF/YV+f93y+YJ0JC5Z30V0Wpvp1IM9H27s4q+bKKdNhg6py/UOXD506PmWCcvkPSgGQ/0zDgLNW1xtAw6glrKbIL6xSzciXb9XYKu+h+7WudMydUoTofay6h2qz1iIvIw5Nlpuwpr7vk5rljwu4NHPU7nU2b2HFxk9Z/GCa6exW9ynqznGoVUuoCziKxy1XhFNMG4YfFfeVe3OPZOV+OpAbQZ/5/kqK42DG6ZSocfccw6BcmhvrHLLcFSb+g7rDKTGNbIhG776u8mPPBWFJZhSdDNs88+0qtEkbUxgPLCGicjt0AyLzRU4F3XEJevCatA8PqOh7h2J+XfHE9f1Ld/LJWilTcfjIYfzamdsRAZFiBmzkcGYo2XJXCfNRBh7xFyNW1qHkLAnMTCkE9moYpfWVOKuUtDfFzJxbxciyH3syo/XUdEa7ijV5c25VNWApNxf723KYJuVr0Jq/J2HxTgIdBfqYkpomA2lj6W/q9i3yTsds912agC3gGOnLlovMwsORB1Eg2XPcsphhGBnlES4y1oT6R6Gy8/RIa4HDwHAGHS0vsTJ9moh3hgH79oJ/v3hGam9juLhsAc8W/7Q9wIhEEJZiGjbIKJymkfuSZ4SlS/U8cRhe/AH8SWG4N/QB7qM5lxQ1RGLs8ata9GbWXXbmIFcF8bQpTHzVqa5af/b00kM08IeACuLi66NMmPfvxsDfcFQKO/053XudfW9k57i3J71xs4bUvIfyWSNmMaBVV9U9ZAGvy79L4kxT9SGyMCq5AjAdTr/kwEDERzu4uYz3prtNWHKYn2JS69VL8ShNufkwBdE9Eh3/g7TubXeZeCUd6/kRTwZVx+WcFoHOchaVMi2IRJyu1ZP56neIXFXRF2ApeE9Dt+lPkfQuiFDPesUKQy47Gjo7L2xYvM2YqBHLy7elJYJuHQaA7z/FQp8LG/ntSMxAIqkAr2PXRGTrbS9B+Bqj1EasEf6+32MnCtXT/7K6wvcc5P50rwLzQmp3Pegam8TL3JH1bFd1R3oZ8Hqzr2gYFHbOFDB1nifTc+9qPQoPtmIvxepmxI8L1WORXYLoci8XjiGFYW5vZjH2/HALwyMFjzBuZH/Ptx0MzUSbfZLjvHkAbgJhcgWT7Z7l+U6zNHLDTd5IsDhJ875ArIH56BwLkVHgUqlTVKN1ujNH8rPY2yG3geI8N09ACcq9XutqvOUodLCCx6Pxy1nJG/By1vUuzBtcNA7VU+O5nOsBi7z4NxG55uhaMAoJBQl49uSdol0hp69Nik5xxO+J3SOJ1wB6OFApQgelk8Lznsdh+XL4kP0zNCB8nr1jA7cqhhyloa/A5aV69Y6bEKSY/YcWBjHrZBtHQBWOwCnAY7s5LoektsvqknB1GIIgSGvbjSbGtZTQhrDnFb3JqHTHeiAb5sNQHsLPeNQyjgwsYweMVhBmUenJ8Okq9KEKT6Jx+jSeo/9XVN2BYrHUueCyOrV77yrlBMVSwI0Tzqz+lPE/NQZKzT6Lw0bCovwwjyGnk+EMakH4Ki8glqI0nBZRgzmdIKWUsAZypnAG5NKSmCo0cadgNDBk+TWERCfdoR25E9CoYroF6j1QhwDbM7ibM8YD5YBwQjCiggabRjqhtKYZtLLh9lNRl+zzyGjundNNlzr5KJujo1/QwJJg4rlSqxz2JBdmoRKorSWga/eaIBsuz+78mUf8vXn6TkoTJv9Z1tYU6isXotaLypUBeMpAwgdFpVEHe4L8DCa/VzViAv3Az6pH6mOXMErGw3zw2KrDzithZj3mG/8do/IX2Tzp/mbLllj219eu7oGivV6xsU6u0phrUrJXiBSHCjUtW77fpugbS3Q8D4trXdsCXiy1WCPmWMZ3zYOQCVHaSWUdpeGNoWcE0voV8N/lBSflr/bAoS0x7hVO26yeweMgPU1Jj5NkokQV0rYpHldbTtsuZAmo5bGNA7anp5/xMAqk+G0tyNiJO8Gme2NAgMZL+VJJgvl1Y0qlb/aYBx9Q4NhGPUORc5v2vhDD5k52ljdOAa1LmFCA2x4GPtQ5i4H+sbuzhhuIiIGhhJzz+/o+rUj4f1+CJ8YRaCIgmeEdqoVu5+lb4hPogPDyswLcxzdQdjlL6+Ty2zrbAP15dA2HgqBdGg9e1RlLSMOqJLTowGGh5/gthdOKTUm8FaeRQTm8Y0gssVLtbmhZIT1/nUFa6h+D6sB/XeUW/t7NxIDxvyE9MQydbCyLC5ScT7FBQn9QeT5BIPU9S4kea800ckej2/aftb1LfdG7wdoHH/tyVrdtyRU7BZtxGSqF6PXEwiW8cOVmieJPzm1iEOppQ52kAPiv28thSUFrBJaY2TS3GT4Xcd0W78Yt32XDTvdKXVHC/21stgkrXlIyIarELCzRCPrVJdsi7x0PtY9lRE6mT/6m37mX63xQ586P7t5XpNLuOc0t4jd8tM+BJ5fwIclfOGLUxU5NCqfhuRaMCNB6IF5WxWysK6PjQJqf1dglx/dKJT5woiJdepS3q4efHS09DP4PToiiQVORySjiVx7wZ2ry9ty4hej7Kcf/h7+2B/5nfjlX/x/8Te/pJ4RN69eHSkaIpJJc9a5Fa8Av1OH2M/fcxzEe4Sjb6eLib/3H/w78ZO/Dvjf/6+/3tErdQWC0QYqO/L6xi/YteSlMiijEKeMa+3ngT/yT/w0xg9+GX/tb1Cz4lGEv+2nfit+7rd/D//LX/l/EBj4fT/72/Aj+Sv4pV8m8XjXw9xTF5T3xHeRbrLa2ozq/U+9z3s7PFcJoDzb6loYyUqXASFhk+M+rB5haGR516jY/k1iNve0rr2G3BBwUPRHI26/M528m9xU5SsdaO1z6y9Q3b+S17u+SxUYqYJR1XsWKl/bli3J7oN/019YqerU0Gi8G0Xh0QPbJlvlHBINnn/9Y0SMcoRwIwo3zDoBweaSUad1/4yCYT6iNsy14IapA6cMMRc/VEnQIbKeQiiBuZi4gAiM8RTv4UEdzhet3zhawTliX7Iy5ydWRTBvz3boMwbGIIloHoX53/7uPVrtlkf2947b3/Hff+p3/V34F/7Z34Wf/z2/kX+XJruur52aDaV2X0V5NiZCz+pKCgQ33cT06HcfY69X/1w88Lt/72/HH/z7/naum/LOOd8wxpNrooZBrvdjr3lzKQ/M+Un7Nvm78436meMTfu4f/Rn8xG/6IZh34vo/8eO//cfx87/vt/Lz5xv+wB/8nfi9f/eP8mfgygrEaT1hoZPXr3JpnQBomC1r/0/87D/2u/EP/cT3YJ7AJV5O4FK5/s47aH3ZaGWSfd6cKvaha74FclhWJGvd5bBHPBDjibjba9sjtB8PmGfj2uodZPP8Pe6Jm8D87xyCw+8Z/p3+Pcu1zZM89ZnPTkeIRriPQ9mAZ7LslNr/pwrJnWvS2aYgbYOA7YhOZF51AKg+II6GALtE6Ubga9FGBSsFAfV8jP5wj8FDJUttJdb5q1xKWxMWxViS6tp8gTJuQmLyJ8rVW8bLKUpU76E3jJFFULcoYS1DOR5L9ODaWy5nZ8gP8aNqShO2caEho8tT8uoR+Mf/kZ/En//zfxn/8M/9FP70f/aL+PCb3srBIjV4wMyso+D7UcmDsIw1hjkCcxHXLQVxNcC8izoR68Kf+VP/KZvsqr7uVRDCsEalc2EA1sdA5dL0TfL+XgSyTox67rUoj+en2CdkJzScC//mv/Eftro0gvM53EYQKBFtRlyPtjly1VvBOeaBn/sDP4H/7pf+ck8SB7iGhOfZqfIqdaB6cFFzLdWHvlMCD7o1ipYTD8188AQ4pj+7fN5aHQD3IdT7z81XmQ9zrV88TgkRxGzE0VBf/3Q6abQjROqgtw+wBGKdcrL6ZVpgK4OXvltdvlrDMZ6N5AW5gLgVIhB6mx2cj8wzIi8aSVhcI8GNI9c4sBqy8evIH4jMKWBI7ETllxYnOUXaKr/hjkflfvZ8qZuy7Azs1SwXRhViKu9y/uWqiC/ECU9A4mwIbhab4ebjm95YG3W5w6dzRPTnu8bd/SIyFueyPRw1Jv6W3/Jb8A/86Ik//u/8JfyWP/HP4Pf81u/gv/mr31fEC/ypP/PH8F/82b+IP/iHfxo/8WM/hB/88q/gF/7Mf4X1G34z/sV/+u/B3/rDb/jF/+OX8Cf/1H+Jv/LXCLF/5vf/DvzzP/+T+LEf+QZzFP77v/C/4t/+9/4Svn9O/NF/+efwT/70j8oRA7/+138X//Gf+6/xC//JX8U/98f/MH78//7f8K//uf8Z4/GGX/h3/yj+/V/4C/hDP/8z+Ikf+x7y9QX/0X/wF/Fn//O/gozAd374u/hX/qWfxU/9Hd/DeD7xG37kG5zvL/zF//Z/xJ/40/8Djc4lvC5RB5wKrnUBcH+EUr76/8l606hNr6tKbJ/7PO/31aDZsgZL2MiW8YixsQWYJmAbGwdCNw2rmRroNDFNAnSTgdWMPbBYLFgk0ElDd5MwNGFBJwQHwmSCVxtPgMFuy5Ydy7KFBiNLJZWGqpJKqu97h+ee/Dh7n3Nfu7xsS1X1ve/z3HvuOfvss8+5wA/+5Dfj4p++E//unWdw+rpr8W9/8g34lV+9Hf/g278Ez7nmJC4+dg6/+Et/ivfe+QTcOz7/i16G7/u2L8SNVx/C3HH3R+/BT//K7fiH/81X4bWfdwVe8f1/G9901PH23343/v1//Gvc/ILn4Pu+80vxss+5HLv1Gn/8h7fj1//oLhwva3z51/9neOO1l/CuByd837e+Eu3CGXzr9/8BNjYHr+F1K5psMG5RD0m7VK8KarIXBQdJuTvTCo1r0IyOvIhoJIqdcy46O0Q7p5urL0hpiUcP07KsM/3VZcgwq8CTTpVEtWnsg/inXY7sU7BOZS44LlD8nQR5UwPSeZSTAHk3wDA3mz08jQRKfO7B4ydCGLx+EnNkoxsabIpqh4lUtEHExDKXM0WJtGEpiMXvbpix9ONIGUTucIaBcsqxtCvlH8T+OjBNKyzLJkpUXOyG8K4A2G09D2STNnRGXsHYx3kTURqF18i4ZguaNbz+dS/E3bffg/sfehLveP8ZfM0bX4y/uPfD4NU9ODx1Ob7rGz8fP/Vv3oMHzh3hK//Ol+Bf/tjfxcc+ch9+/Cd+D8d2iO/+3q/CP/77r8AP/Ovb0R249ORF/Oa/fyfuP3uMk1ddgf/xJ/4Ovvqj9+H//qsn8Du/9g780X+INORzXvoC/Nx/94X4iw8+jGYTDg5mHMwliT95+kp8z7e8DD/7v70Tn3p8i1te/nz8xH/95bjzzgfxoQcXfMs/fBNu2jyE7/+Rd2CLCW/5x1+NW44ews/+xl0AJjRDVii0P1decRluuO4qjBWPq04fAKBeAhMODlc4WB1gaivM8wGuvPY6vOVrX4Cf+Z/ehvNrx5e8/lX4Fz/6tfi+H/hd3P/0jB/+ga/A7/zPf4A/u/sCVoeHuOWmK/HM0Q6//Mvvxgtf9K14z6/+Cd72kSexWW9w2bNvxk/+yJvxgT98H/6Xf/UArnrOTfjn/8OX48nHn8Rv//kDmFcrfOGXfgGuvPsB/PiP/z7OP32EXQsnlDfeqeTZ6g4TDFDfpkB1GkRtakhUtM/J2i1To6h8UgENNoKxrT/FVbTjlmihlTOAV2AEKCXw/GyVyhf6CyMhWy0Em/y5nkSm7BXZLAanNmZasYRPflI8klD/HOIypXYxsJeQIyCO9PMk06T6iopOei7dyq3ovSeLhsUIMkmJoRp2g+ZuBjza5N+P6wdQCIMCIrCkV1WQWKAitoCckG1yGlGdiKY5bpravJmuwGIyNsNFeWTlzYLVXQw5C5dLyOKtBXfTTs5485c9F7//r96LZVnwjnd+Am/551+MZ/367Tj7zA7WQun5nv94Oz74iYcBd7zjTz+Of/A1t+Ctv/0+3PvpC2jTId723nvwz77qWqywxdpXuOuOv2ZUaPBHz+H9H38cN990FfryMDZLw2a9wYnLr8Y/+vZX4w9/892488wlSBSmzDTSFeDtf/R+/NXHzmCaT+LR93wM937Hq/HCG6/Ehz59Hs9/4bX40H94H849FeTYez/8EN74+itw6Wib0FpcViOU/q7veTO+k6MI9WuaG878p0/Alx3apNkaQHEEHb/7ux/AJx+4AGsT/uD/ei/e9JXfjTe8+lr86ruewGSGZsCFC2ssfoxHzl6EoaEf7bB0x/GlIzz9TJB/X3TbrTh1/mH8xtvuwTPbLR4/fz/+5P0vwZu//Fa89c8/DXfgypMLfvYX3oMzz3B/c4Ypn4l8nEY8Giw1F2o91wi7jKzqSMVQobCYzjYkUclTTdNhdPeC3ICDzgCJEPYnxIXuI2ewQim9Uf1qaZbibNq0qlS5S9YuMV21W4y33SUa8Tm5oonIKt4VXBtN5KLUoS+u21qQuX/fhYgpczZkvh0HUdOIUFCLoh7vnNGwbPLhdaN3MvygRBlj7izkMGs1yhJJVkmCHd4+0o82naAXD7gmAU9r1XjU+w7T6vTwPfGeeTs7ndA0HWLBBr6sWS4GdC2ckEVOUOLz3voFL8Irrm944qu/FK95czhOXH0t3vya6/Eb7zmT73XmgSeTc9jtOtbrHZ54LLpwzSasd4658Va33vDClzwP//nrbsVNzz6N1QTccutVeN/dK0w5t7PhG7/jK3DV43+DX/nj+wGoaaolLyFH/OCnLpajdcelLXDQAIPj3k8+jtv+1q1420fO4chO4A2vvhl33nMfAmkGOtM8E3nXn/vpt+L3/vIsTDmvAW/6ljfguz4PTEWk5LQ07L7tePjBi/H77DC971NP4OYbr8Xu6EH89M/9BX7gLV+Fr/+mi/iTd9yJt73rU3jyiFcIALlOZhOe9/xn4cZbbsav/eK3yTBx+vJT2N1znDvz+F8/jIcu7kLstmzQbEU7ZmmaXc9N96WoWiIOjgewptlTwKf+CiFtJ7eVXcckIU0NfVQ1O7mdAYkEGtgim7iSv6j0PCegi2ewOS4AUtObRuWRX2g2c0zipUDTSqfJcWmmqgK4nCRI9sdNZ0Q2mLDkZV/BgM5wN5WGYEab2uZBdW5I3JFJQqjxz3xdHpW5ly1Ir+Z9AZYNfDrAwivdAGBZYt6ibu3O8pbyw2XDCcTrdCiRwoCfL2n2MZbxhnU1XmULfDTxgGmRLhTKAbGEXO5xcxqA5EqkqYCr98IT2XiLO1Tf/IYX4EPvuwcfv+/xNLTl8BS+8g2fh996z6exZml42W7TWUVZDFh2a3Te3r2wPLdsL+FzX/n5+Pkf+lL8+q++G7/3O4/g6aM1vveffhPct1h2x3BfcOurXoZvePXl+Gc/9ic42hyjtXDYyxLCoN3m6ZwKvdscY9kdwdsWjiAWe99i2V3Cb/3vb8cX/8w34+d/6iY8s1nwwF8/gJ/9zQ9h2UZJLYbPRNWhTwGZ+3Ic/A9LdIkqncFCPmJZoy+8ud6A1rZsfIu9mKcJ290Gy+4IH/nLO/CPPvwxvPyVz8ff/3u34Wtf/3x8/7/4EzyxkyT8iNL/FXp33PPBj+Of/uLtueetHWDZHOXB6LsgswNZ9tASwKGJUiECbMOzc7iOgmCO3lPz4A6gitF9iSClwTweUn54D4qxL4EKlrivI5DzAiBEWm0+CTg1DEn6tyS3O6r0CqgXK+6o6cbzoFIyACzBZcTNfzNsp4u3HQuO0i6h0i1PgrGcGhwMhzANfiD8pUeM9y36srM5AJIGfszpD+NgSBlGWGsVmeMD1SbLw+gO+JICpWC3VyyBrsOr+1KDRTRyHDXTATCggfdyULLKnG5iKUkcAwBMOIHqgDUKYhrLWTu4T5jmk8PGchJTX/L3O+d5et+h2wbTdCIHkABqX/c0ODPDFdddiS97yZX4mR/5Q3zwgUvQPMxrbjmPX/+pr8RLbrocHz0Ta9CmE5gmGst0ABgwTScwTRtEeTNKavPqNF79qlvxyF33463vuD9MbZ5xzTWX44zHVPPVqcvxg//k9fj9/+Nd+MSjsSbBFQCtRQl1mk8NzW6HmNph9AXA4uBOh5imk7j+eTfj4NEH8L0//R4cbRZsd0HiTnNdiwcz2BTlaINFCdZWcE15ElqEQQ1oYR8hXDI02GrCrS+8Hh985FG4AW11gJe/+Br86bsfhUrB23XHh/7qbnz0jofwq7/xXbjteVfi7fdu4R1YHR7CLHqB7v3ko3j2t30uDrdrPPTUBq1NmGbw+sVCpaLz4MR3g6BNs1J4bgK5DGg2hv2eiOhLW1eLv6TPCevN9m3XQj9S80gtSfhOxDDNJ5GXGQFRJSFCaNZ4fWD8bJ4VNZf1Le01UKaIfZ1dazOMneFagoh5HFOg9zalqoXyAV34bTlYJz5ghk2HPve+s8aykaZnayHLM+7qS6L0kREiF53eFWw6qryJD9KrUQWqlMDijhInHWiWudOyOy7Glj8T8l5km7FKQtlIJcSBjkUty95jMhOoI3HAneKvZcgziZokEopW9WDHkRvLiohNeOVrX4TlwQdwxwPPROOPRcpy/lOfxgce2OLNr70RH33rp5iyb7BsL3HTJJxZoy8L4vqLEhzd/+nHcMubXoQ3ftFNePSo4bVf8TI8/2rgDCX43/yeEhFlAAAgAElEQVRfvg5XX3gY77v7HG664RTgJ3D0zAZPPCU0GPeqej9R76aLeiWw6+EgL7vyNK646jJ84Stuxnrp2K43uO++x/DEUxyN6AsaRxf2zlmpPtxkxf2PjlGpZWlgo/DNgW/4xi/Dhf5BPHKx4/VffRue9eQZvP2Dj+Pw9FX4zm99Ce684yGcf2aHW158C67rT+K+x57Gsul44MHzeOObXoH7Ln4SFy48g4/+5Z345Ne/DD/xw2/C//lHH8OlZYWbnns9nvnUvfjjD5yBu9LpDlhUIHJ+BtQGIH5Now6mRNFBcrJawMMcZl9NYtIuFMTfZYUsWiBC+dn7NgjHgSD2vgsZNSwJ9zxXA/oB5fCgrF3NjSH0itvZjYg/By35wvm0sb/TdAhNvIcZAjd0HqeYMg6PuSMq2Wa5mNxgY8Wz9y1mUHThzlwdu3yoUQ6twSG5OH3DHKqhL8dkgaWWq/owfIPWD/Jw+3j4s87taFNNKvBlG/++bNCsnJGzFuw44IsGF+IkZYp5riE7ncgh0ib2Miht4bWCxnxcU81dY+2oiYeHHiKnOrUZL7zpNN76+/8fFtc05XCv8AX/z+99CN/+xddi5ffinrsewuNP82Y2A5bjNe686wwubZ1GO+HS+afwsXsmdDfc8a478LOXOb7m734RsFnjPe/4EH7qIw/j+e0S2jThhssN5/wE/tvvfV1yFB9510fwy//vvXj4b84Cjz8ZB3h7jE/e+SAuHKkTdQ13w713P4Sz56O0+6zThkvzSXzTN7wSgOHgxCFufvYJ/NS//C28++MXIooZ52Fsj3D3Jx/EY+eeAgkd9L6Gu+PCo+dx1yEVog34m3sewqVzl8JOdmv0zRa/+L++E6/6qtvwX1x/Gmc/fQbf84N/gYcvbNBWGzy5OcA3fMNtOJwbnjj7OH70h38bd565ALMJv/Rv34bv/a/+Ft7yHV+Cd/zBn+Gev3kUP/aDv4mv+7rX4Gv/9qtxMBkeefBx/O5fPom+O8aFs4/j46d0XYKnwldROLaz18FD2N6yOw5kJLsNq2dkdbjVYe9yQLSnuM5imPqm3p9lg86+qib7I/GsJjWQ3JQjm5jixB0nnNiVUgJ2uvYtJjsJoSh4BHSpp8VMSCcTDmiHRm4j0w1SUaoUjVcDWO/REJfq1gZ7+Wu+6wk7eO41cX7VVLXkoYMIs2Rthz4J5jWqFWtaEvIrqyS57NaYVicjyrHiIignx6TN7L7Ln9EluTXbUZqIWmCVvNIbTgeQtFr3SUqDYTDCwGH8HuvYkZLsME0HFH51WC19QreYYnSMmpVAA7CC4+59fwOyYtRqDVlxaNNBRutANcdp3F0SYUM5uSQxgRogqwiqEYat0qxc+w3R6YQX3vYK/ORbbsV//0O/j4efinx1PjjEd/6Tr8MtF+/Cj/7Sx3jjtuIr32mqYbXqjUlVpWu8ogYmNVx+ww34tX/z9/CT3/3z+Mh5EdhlG+47TJP2Y8q1KgzNakIedA2m4d7bjGmOi63yXhir6Wk5NyUncoE/O+7FnIetUnB1QquC0Ya99ixtitgUmt6TH+hQ8n/dO5+1+kBKmMVZK/Mhlu0Rxo5XjWPQPrsvmXqOc1MqGPdK4RXgfZidIQJVfU9CPa52e71HrddydM+FJm+ZXq4v5aVQqrUaMAKonCbYFs+qQ8K6sQM1TKUakqpVfR5yXQ10adykuG1apaSm7tfxP8ZxYMPPx0E+qO9kPtmYR+vgZz4OVTqG33d2b3ocquzcS4m6ccM04owRytWngoSqfW9UPtcIiBxRf8ZDpxQqhT7DfxqH0mpKkiY1679yjPHM4XSj0csL0rpa88PIr7zychw0oKOhTYZ5nnHFNZfjpS+4HJ964OlwYmmggKT1I6M/ju4Xh2E08HzbPRJvSRurtagqQ/UeAVKW9iV6LBb2S3T1ZuRl3dqvnnZcE9O1VqiUtG9z/7PyoP2XPevg6bNN9mZ5oMYhxarWGRWQIcuuMQjJJUjFmvqdWNe0Z2uMSVM1StKWsw2CSANeDiLTKVb5XL0gdNi1H5xYJzvu++lYoZfqN0r/YGxR190UEbEmwANR7M26/AwRlhpPZCRQeYgH3ui5Td4rHUtND/YkgtTnENA8ZckZAYCQhAwzqQYjDGdFAUvfCTgyUvBMKjJ1jaUvYVd3EkYs9RlQhyzbvi2RTR6Cro48cHO0sC1nGQC+7+FZMpPzgMccjEXakTQKSsL7Alh1hEY1kdEWlsIazVzIuE2JsPQxzaZEc963+PCf34G3v/x1+IVf+A4cPbOGTRPmBnzgvXfgN//0oXJC1tPZqneipdGWG1S5fRzLqMivA2DW8wDXNDLC5jZDMy14umHtAG3QBULIUtF8EccmfopO3loiKI0FiKPZIB0BvGf4qXs2+LeGLtWuRxJmp33ANZ+k7CJ7daDb82pKlgLtGNWhEQUZrBxtCASBejRPBflsPdHlikhnx9kehrjEqg3fGe8JyAGjbFb2qvJock50riRrw4l02Etf9R3nMN98tV5S7cM6LAFJaLzDzWGV19lwuHh3BRlkycNjlNwzkY+lx0P+vAi4gFFIJ7LsjpOYiwlSQUZlay+Uq1F3L3nqoPCMUpfujozIo+cQ/BMjDCIppQW1QSuohKi7GZZlM7DLBa2T+Nv7FShEhzWUj0zxYDltWQhGkDy0QL0MUpEto9SSkBiDTS/LEatBM6PxGjMl7/GcEik5TpycsaKQar1eY7sTlxRTnkwj5wZjzdSSwjtJjaMNfRTkATbNOHnCcHxpjQ62ppsQHcVIef2eUt6wIZvmQmBw6hGqR0hweZoOsfRNaoDyu62lDcqRxeFRR/U2gt10SH6gKimpnkwb5loyla3UMRq/+hIT1sO2KsWBlyjKwQHJmMppcXFrPirS+QitL0vcsZqotoeGJNfJDMtyjFSUQrIEtWOwjcGUFle7f++bSFfTcbW0Vy4GDI5lff+FudkKcWP0xJ4IzSXkPZ59W8KcdoDSUNQmGGFWwkIdnbYajGnBNJ1MGLfnbCi4MURw8a75liCPsipCSJarTefPTphzMfN50EP8xnzVu1KIIlbVYdimAy54oBW1n+vrDLyfJI5MdsiOald4QVYdBHAtYcaZCWPaVIig66BAcxb0SwhNULLWLOB6pTqtKfdu+Q4qCydysuJMAGB97Fg7h6jwkusk+eYT+w647+KCaY6cb9GwTGQ58AtTEYpmE46OjmB2AlOSgio7eh7iuGiIZfWhHI955Gnivg8R2VIc692sAXnpMgNLm1kFakQXyV2wWdE7WjvE4keY2yEXWLn8FPNMhfQ85o+o+xMwHv79IcGaZ+GM8mMgiyKCTkjxfuPl2QoW4r3Eq8V0sg168umqNjFV4fStcmJKnzlzBpqWVWrrKIXHnSh5ARVCY8Iv4f85IkxwXqRz4IWqCdCEIuUx2QVaET0bWrpuRWJ0pDMIDcVhVB6a8sa+t4DxguwYFSSTKs7DazeMB4ibpFkCxglHxkjEP4ucd5vQONOe5C9IbC5bdITSb8FYPYmGoHSQhH7G5+vQbVGq47T6uVxo5Yb6LR8iMclhRUsSxMnMi9eRGtamKBXLyLzmYehzRiOKvYtcVFPUYwhOz4OSOTjXI1CW2sC3bOBjExRTi3i/asZyGrwQoPNn2zTDsRR6Y8QFnZNataMfB8xs+Of5XlT/ZoApuBwpp8E1VYr7He8WupO8g6NRbp1tAQW3HRMaNC3LUAQ07dqUOluWQTWHovPsyA7MioQPR9CjbaCpMtPSYYcdc+AwwnmGD+l5V64j7gqxOeTpKUugfEEpde8bLH2NaT6BZnMEPlfodqAjnYzSneSFXFPnNSVO/xx/NxZs8tl9Z+YLMwcRabth4+lptJl7FYLI24ND2CHIqoWejKkJmDP5AujiGzgbvHouZjOO+6LhQzXjZQ3j308CSo0z+Vn8rhbOQI1sDmBqK6BH0073OAih01inOKcUmgvLSFHm7EsfIGnkmHlPB3o+c6UeagGXwTgKbg8CN6jS0WH8O2Lx4Z03gzFWeXl2M62bhfaD6Kolm87PjRgCONeVegO4RxORIkiW0DpCJ8HavYk38CRVNZEaVrd25whAm3KUobgKIAbFaAQgj346p3CqvF29zdW+3caDJwWlfo7knip2fQdrB8ghNj2uf0CnaydvFNTIMrSmjwFPzjXGF4Tj9OKYFAhsSqWmJsdpv2xYf72XoYY1x6Ahnhvv+TMiFWUVzh4QQEWC2LPW5vQj4qOEcMG1DiTJcivXWKgk0lXZ66iBCptNvmmPHyHqNssvnpPY6Z3NKlwAQTHUL6NXgrX8Z3mueEWmGMx9VMrJiolVZBplqHH+S6+wn7MpAg7ir/DJELGVV/xxIzDUxIGhSxVWJcom8olOL6PmyKqPhl2/11wpADUIQ2ObtUERZ8YoaXz3OKQaex/fZTAexC7Ek9GqZ7oHGHwZnRErSLk2lmRoQPQqP3pf0FaHwFJIyNLpi6WUcUjPoj0BwAE8YwqayEwNT8DQR9J583tFPzm8zOEJdXXLvI1zUqEKmqIrt95a2BgapAeKdwl4vWC771TANddcVQVJl25G36YICtqPnIBQQM+Urt5Fgq+yBcOMRmS9bz+RErkmljk4T1brQbJeJWj1fAyBAfPQckAnXvtnuQdCRFEoGN4fw2Qx7+zPKslDzCcBcvxD9pzE9/W+tTlYWwmZlGrQULmxbeLLsxM0eiwKBcTBiHmAPSH3UDZ0aikWLqQBPnhA7x1Lr3wwDrQujSm4uKdrkA7E82XK0BsbymzCsqyZpmA/+ubGezqJ0cjAPDFSlpbPJQMtw0M2JIXh8ZAyv9XVjukwOdl8bx4oCo1EZ6MzmqsyUsgkZcWChwkTAd2rWurKcHIpQPNw4k0GlceQhOeg/Ui1oiaRu1GDosM2XBQ8lUONq0BplB2QKrcvO0zzwZ7Tt14TukWwOTRTpZ4DQmxdVYaqhEllON5lU5dJx4TqsAnjHvjwfrpTFLWuQg/8/iSlWc1IIlJdqX0B2MAYFbAaIpVj8noM6tEMmExxVAkCdRrsuRLi0D67I9Sc+jnZJuQs+/6z6dC70FzYubRKCoxlk0w9MxWqEqvAgrtjbiRv5KAUySOfUo/HAB9V6hlY/7pVemKeE7A2PGrLFKe1Q+hWLxlokKkicRCGAeXrO+gKgipnVYlLRgR+flwBIEJQZb4Yl5Z8iNKqwSvHNYBLvrdKkCrnKidU3ToG/MTMz85cFKnPr8WVAm4fWZUMvQQwEhxJNq3gxlKXRZt8pTsiODvVq8hc3IxTyqgx6TuHQdc8jOP0S18CDORpkouasxBOKN671K8SkNnedQIc+dYK6uvnI+AMzVsqw+Zk7V7r0HcQZxODxHrunZmIPrZU52hBXidIgjlLznzG0tPIfhuqbZ1R3WQXSDvIngu0SMGGQc+kCCEOYtI9NEkgsk+JKE0p3F6pW+V1Ip9AMEYFZ+cazBBnMk0HQeFA6bECjcE4WrIkCYOT4Lkr0l0O2tCmE1h2R2zgjInwHh+0h+TncAozkDXjyI2dkb41RtYcGBI3TLlPqX2P9VUqIsewSrFSS4ZYyjcg7zdg+apEKSqPKkKjNiwlslWuVPRv1hDkFNJg6hp5iXSGA2o12CQiphwZiTx5/jYhW5EJgfPSYSC9t8RFKtPW9CTmxpqJiIDefSEcb7WBeXcGD1QzEGWkCxqcKh1ZwmI6ek1/akWMpmF4GG2zFVZXXIbtUxfTGDAcSB1wM763KZeP75kODuG7qFx0Iih4h0YE5DgBi1F23deo9v4GH3Nj9/BzUzVMAauMrK2puuGY5kPsdkc8VOxCZlUKrNbV7zek6hIF8bVcrR3k9Ku8TS3+IiF+YxDhnbDkvALphn3VrV7qpvW0a6UwSmMygLkQT6k/h12MvwfOvBVxKi4GU9kKrT/XVE5gikl1gfax92yV7hQRP7ZGlEKYTrIRRJBYbmo6cUJFwbPIxWMSc+8b9o9EzT6avKq3X3BMI+vhum9xl15WLO54x4KmTovccX5GliFFlA09KbkpgxgrnwG1kZqFoMXMxVVZLX9f5OoybGSnNycMhDysog0vnUGJb7IcpuoRGXyDSoglttHPyHjymaQ/cOfAXYqfQKihzw/cDM0QkWGfeu7z8OzbXoNrX/kyrE5FiU7RK4a/huPCdIDrXvMy+oi6DwYO9lQt6L7gihfeIowFa7EODuDZr70NoDRe079liKqUqEQdXZqeRiuhme6VydRO/75sME7DXpYjtrpvQrgGEYOyxw2rBBt0590hfQtd1qx7P7OS0DvHGKzZgq8mxHh2Z1t78lG01z6QwdI69L5O26zCwJJ/nu8NIPtCvOy5AmKlkkhnYMOfoVAlnW6h07KRIlqltwBLuwNPJJRLh5DrSYcG8WbuqXEhOva5tdmtHURUM3mraBtPCbVpiIbKd8r3g2QMGCqFJZD9CgiDiYeK9Zg4PQoAL4+Rt7PUFzgqDZKUWLAt8raQnyqFsqbbn4prUIXMB6cwlgUl2e3LBqFCVVfmgjadzMEksaw1cwMeF8sGcx3vFocfUL19VItC/qzX2qhxLQxhAewAams2q1pTPOuGnxt2oqEmhkJGzWZc8aovweH2LM7d9Um0U6exOnESy9ERzXjh0BmivstvQL/wGN+PkRDA6prn4LKrdjh/71m0tsLq5AmYrXDi5hfg1O5xXHj4AtrhtVhhjaABGtwjt5WNtHaAZRdVnpHLUUUpxdUiv5UuBsgdHCzXSlE/06xVRs1AUAdhU64AwiNhjWXoUQcUvIGqfOoJUoAzouRcV0RZFsN9snG51kEKvHRYUwVsQbYmpxObD4kWU/0qO3ehqfre+Fy+f4tb5WT7KmFnCuRxDhYGXoh3y5RmCwNTMdd/K6DHjBnLYpcCzKhUlkOdrrv+FT8EnD7ZstYeeZ0EL8rtBS/d2UHpJWoCpDLU35ONOETgwB3TFN2iNnhaeS4wfdAt1fqu8nTjZTFi2dPtxCHPy2tqzH8QaFM+V1ZPgGo9T4TiiSr0z57f23MNpiYBUagYW6ZHIhot/1//6Z1TpxKOc3fMynnAAE2Hgs4Dy2fsdUmSlt8nRvtZX/QiPPre27Fsd9hePI/tpWOcev5LMS8XsVsH0XbVK16O9dmzOHnrizEdP4nTn/dSXHnrc7F74jG0y67Dc77yy3F4+hANW+z6Iab+NOz0Dbjp9a/FdLACdk+jn342DvoTuPTo02inr8R1t30hrnr+52J37jEsazZyoUMKxURnXaMYhQyBspVyKMXzjHtLiG0SRpHoFQJsE/pynHuSa9fjfpac+C4nNVQSxpZzeU1TSoIxLbOyDa8ongQssPf5Iy+V6lwv5AsgS9g5uo7Pn4JBM15atU3bAwdkK9Uu0rsOulLVVDq7LiUSIgamJiK5D2ssDyCHIRpgQl/OHzezugNxlC7Xyw2bBgqfxhwsfzXqAz770ORi+vj/Vp/lijQ9FxjMsRqJndwkaE+12TseNslUKQrrnPI0CKQS/gnG8llS8afcrsccRc0CiFbr40yrekLoMNhlOab4RxfqBLyO/66zLLUIMhMSx9yJz7iEBiEs8r4LOTUd2bIcBSfCIcNVfg3Yf3R2g6teeCPgBe0vf/71WDabgL7TKVx+wykADaduuBYnb3oOnvzIh/DEx8/g2te8FNtzZ7A+dw6PvOfPceHeh3Bww02wZYPjh+/H+uxZnP2Lv8LFh87j9A3X4dJD59BOXokbv/RVOHf7+3HunrO46sXPSSNPSAtABJ5IOvUg9K6yNY0SXvoYVlkqGKk7cyS3B5gu9GqSqsvBTvkM+1Lqiu4izuNmeN1zQttPrqic/14VgdF7XyIgYjei+6g+HeXYdTgtbVDFhdTc0GbG9Ds+sxrvxO2kDEHpHkuiy7LeS43KLpf6eQ/Zd4wcCLvuTOWikrWG911rWVLzulAkPGNP3iEerFSaOlwjbxHj1pZhgT1foGcnG0urZtB1iYJGYw5WNzch88DiU3bDz4RRpvCl92zP1uU9kUv2YePA9MpyClKzacjfgMYLh5q6/WApGW9UVba2ygtus0OQnwdGgeAqeNkMxHW0RBuNF9dkhyJ/Jqcj2UwjjOdTypORI2Oz4cIH/grLietw85tfhxOnTwCYsDLDdh37uXr2Tdg+dhawGaeuvxxPfPAObJ5ZY3PhUfh8EsABVgfH2B7HAT35rMtwdP5JAIewdhG7zYK+2+HwtOP46TUue/HLsL7vE5ivvg5Xv/hz8PT9Dw8RNW6T6+S+lmWTxiu7MNTtZN47DTNsS7aiQxRIc4LuD+2DDQQ3MXAB/B5nyuHLLlCHbq9noEBfsIcAMJGb26RdCc7L3rvs3nXDV6ONDjeWZaRWyRnwLq7uMzs7xfP0/Jy9c6VAJmeA0uoEz0I7TrpgylRePJa6VSNVi6AsW1d3si7xUutDofmwwdAxNW8peXEZ64AWMkqkeYcRSxorL88BvBhq1+ndvLoxa8GWwRHx8ALDwg+zEWkQaTg+PNewmPDSWlQVxAY0sEuDzSvo0rsuSeBqsI8v2zTgMBh9f2xwIA8StTwMqcsg9EzDEEzskiuDB2RTCEUG0Ts00i/VdwNZB5fmYGjT7h19d4QLd3wIZ973Cdz4FbehrU7D/SKWbbzr6ec9B5ceeBA4OAV//AyePv8UfNliOnEl/Og8cOoK9CfPcR2A1ckDbC8taFfdiOXRB6GBss0Mu80Op2+6DtOV1+Hw1IzH/uzduHj2qTwo9Z6s/owHYWjbl05ijIjote8ZLeXoGZgSLHcRcEIYRAAmFCrNitWz6ECkjfeK6B7PpMoZBM8z1/dAh0SzOaM0S8FEHHp/fj6GfZW+xbzSmJycjzGFCd1EY5UtCg5bZOm9O9Hzvj3rAvMgX+uKSpVJJf9PfRPnpMa7lCMXMtQzu3cO7FVvSHY7MkenxgGDd3OKtvKlm6Hq9lofMcDVMTlCJWn8JTTqvGs00Qahafy8p9cOZ7VASU55mPis7IRsVXsGRg6B/yvOowX30lm6DQWs5YE0F4/j2eAk1ltwUlcvAlK+RX5csx5I/pI4azZjwUJtyVAiBnKgiuZ5ZPu2VYoV694RNXWHBHS6pbtfugRME+zy67E8/miswXwK1770OnzqA1vM116DNh0FaoHjqs9/CZ6++/04uOZGbJ44G0s6ncLsF9EX4LKbrsPRQ/8p3uXgSmD9eKC8ZYPzd9yOo+MNG8GI4NrgwNEzBYN7zHDN3owl99/zwHquRSgQUXdw0nBJKiA5HlWf0lGFA5GuRvfTOKRYFKncEplkB69LByFOo5CCM+XTHnXNxaDNaJiSbC4DBPsksgXckFPjtH+jxkhBTt2hCnLNDiCeK+0B02AfrHpZQy6ZSFuOOgw0O8NdVTQ514nK8aUQMc9JUE+GZnOfLYS5cVbz/kZ59qp6xEJrzDuSBNQDpJiLrG98h0GDQVzIxMC/GzMunAdrrHqA3q0lCxzOI8mfFJzIjjxzz7wHVNcZoFSnIlHB3BjsKlVqMKYQItLiveszponpgG8xRp9sZ9YvLwGODGC8yd1RgquWm73wLElroYMVa5q5Lkk8ZXxXv/I22O5pLDvg9C234MKH/xy+OY3Vsz4Xp56zxqnnPRf+2Fksu47Tz7oGNl+Bq190K6arrsd06QGce+QiVjdfjxM3PheXP+lY96uxO/8oYIa+2eD0LS/Btp/B9sTN2D72CJo1XLz3DG544+tw/q8fxOrkChc+djfQZo5a5EBfOtKOMdIabWAu428ci597TEcBMv2+Dkm3RIJmiGHRSulaornGK/3iwEuJGRMsw4FH82HY7jikZqaeJOZuxC+RkRK0NSzLMaQjSjuKaIaprbKBslG5ObVVXAXKtw0Ojg5JJXeeN1BdjPEctBnunEuiAAsFZjqbXpO3hGy1NvHNE6eeFTKPiXYLfUrPzzA4HXXI6JNLBDBdf/0X/JDZ5SdVgtsrm0BEZI34GqXJKgdmZKXBN4suPh0KHb6JhhDuyWuDqZ5rJClBlBBIx+q2JKAcxtinIFUgSR/9e6kFSU4xUmcPA4amLBgh5S4NVrlbss78MwOiw4/DTWrzgrFvQ6QSIQ1ElAzxy5ToyxRtpBB1xPUGqAgnwk2OR5xG+KQddk89jbaKhqonP/ZhPP3oeWD9NI4v7rA6NFy8+y4889Dj2B5dAo4v4cm77sF06jKsH/kbXLjn0wCA5alz2G0nYHOM3dNP4ejsY+ibXVQ5bIYfHWF38QKOHz+HvnRsHjuD9ZM7TFPH8ZlHsGxqBF/nOiGd7Q4i0tW8VirIhqzu5O8ztFgFIdmhuB8hreCW1P0adtNItqv/R52eTWliU1vBrr6bz5rDmkw8ldIp1D8PLQPR5CWCcmZkJ0kZG0RkUIpLlcgrkCDXpTprRfZLAzSoi/uOfFmRtoCnrSudtiy1IoO6kH3OaPFosqz7avWMUphS9r6cW8/lGBe4S/atPoAD3rvITXQyHCIKvYfPHrpMxU9gOEDRndrhxhuQJrLWXRAtuj1TMabmJBeUXRI5SHgjaXkuKo2pm3JmIglURBabjS5HQk4BAU2b9CWZ51J4JGjpHY4tnOVOQdFS1TnnUshhiUehwpGs/x4RZi06ElVy08xHdyIvx/hLCtKRhV8uPY1nPvUMlj40CqFjffYhrEFyenMRcGB94TEAjov33Vt7RkT1zAP352HNqsJujafvu5eDftSnESnW+uyDuNSVhlBiPZEzanT4GlJj4o/o8BAooXt1D4cN2l77vIMiPqeleg99Dm126QswnaiD2XcAn89zLsQSfJrAqPJypq+a/m2w6H7VeUCJCutQxz0kRgK0SFtGZLe0t3Ag0dnctZ4KRJlSzGlHUteWPiMqZGNA1t+rzlM9k+bYlrPNfKQv1AbJgYho1QBh9T0pVYqzOjoX98Ub3E1oYVThhQcr+W75frkXvUBF3yeIU9wAACAASURBVEAILeFZ1H0RENoqNxP/ULLTalqrslSVScUQVxWAHlWiJ0YMETVyNFVGKyGVHIYIH31JsxXJHF4ZMOSHKc6yQj56bz2fHKh4EcHqSh1ULhu7a5l3yhDSUYhxpwPKJinl5OpslZPZ0sgVfWvOYrLyGTFqzffeR2s/rG/e/YKx8Y0VAK6p3jhREISs9C5ycJvcXxF5hQyq+iMorUMQdrIqu7JCFgWdYy2bVcNXBodB5l6/8gv2RFLg+kH9JRnNFXTGj9gXaRuAukTJcu31DvE6KnUi33NEvgEodkVc8vuL4Bc/oyqLvk/vorkeNUcz0ntPW1TDmOxfvF2uFcRV0LmDqbt2oEsy7GUsVesGypnoMEc+U8wpqqvRVWPXYhaEjoMxp1eGiERtkgN7JFcauEqT5aSCoVVnnZa7mqWqmad4iNHJ7TslpS08uMnAC+oyPeP7KD8sYnOu0lPW6ie2XYfhTXYA8CBV+YoTrUxpUTQK5WBcpYE5jUml14LmYJkvdQZ9GLUnOEwE4mxLRpbdkJ83Rs7a9ymfv0pqJZ2fbMVysP5uvIbKvPsRdKImMjiAqnTIqaEcmJfatJyG+CbUu3yG7fQe6DAdKVoShUop9c+17zpUYW9VztcBLnvUuoh3ACwrKIDhs+eQiF9TGnCAPUk1z5K+Q58jzi0cwv58k32eRuvDNFvOFY1prOfvVUpX3d06AyK7p3YINSLmuRv+zuyCu6hKR6ymYJpaa7nUXb0e1PQzZch7FbVIqCqItXIQeehoZDkC3nt2mAJIEjHDk1saSzoik70NUmZTbTjGmekMFHFaKraMALkVE9zXJOmc+0gomDwI40xGTz1XleZiwyOFalm1kBMuBJfcxtLZtKT0x6IRysUB1YHXd0fOLYfY6llgwRfJYaEIunTQ/NwAFg6YDk6kRTqA2TjnO0ytoSunpcU4UUkgyDD6Zg07OupqtBommRM1aRRe3hYjUh3U4QhJKVICUIerKgvuHR07NIv+lEiLAbXlq0HROXmqgZyZBZme8uqUYxs02BhKLaSabTrMshYdWNkQHYwyFgcMM/LOUDN072hWKMLG1XTERC5E1S0k43EWY58p2oKnE0c66Q51gTfEkO2OjplNeCq3Fg8hW5ny3c3ZMJjBYMgGbMYC99msmURMOepOuVF6K4NDHk3R3+tLk2BEOgjBbW1KOKWY7JR3GyQxxLRlSIUWrOlIouoS2nt5f4d4i5wp4A40lBNj/0jvO8yc4xj/rZkUKq/JCaZcti9Z7VCLO/jedRuXp3evQcalS8nUA0v+LP9Gfj/g1RegUnSqDks9W0NiV4gLbYDWRJLJmVLabhOl5QfhFEieTuyp0F6FYx65JkVPpBMYc+kUTKFBUm64bCYIxN632O3i0h0zFZssD6LWOPZhaETkPiWi9FFs5zwERCSZmxepHn+nGqZEdnobKgV7ZDt7TXqnBEOSa0CXYes+EXPOu0h0zPewzmlriuCOnlxVSQZynogHYsop3PB8Z8nYsXRofssCkfix9vOkKzjH29djZaIjPMyte913IxWm0KQcXTgPKWIDsaVsPOALxkxC51czwFOqrUGlgnYapzemF43RRjr+7srzURBGm53NW0uiiTDMGY5dXFCrkipZ66qYtPT0c4u7JhsaOpZMZ6RLUHNbsxjxVvc6VElThpufIfSkyC/kYxbOmn+eug1Ypj3S2osT0bOgDxHAE9ymIafSkwcSvdrm+cGx5s5yaf6M53SjBjH2EytFgppS8nEMG597YkRVNaAxNdQ+av2FDBgKcj1B46/I2jI6mzdMtuIdtlGJCGQQISZ/eZUD0wGnXVlWimp6WR3sWC1VUQQnlV50Rv1AyJVG6tZwHV72M+VnVFoSTYRyZOLKdIh1aKs6YE47NMJ9cyKfsWpoaodMp6bz0iCUMeWfN6E/OXMG6MaKjg63Ic5kTjnM9ehw136B6x97LY1JUgj8TwV2z0bDmnSvRju5GIrtS17KF3BjtK5hrskNKA8aYKKRCU4BTeajneo0avXFVXD7dYAVGcFDUkRmPEcSYlqgOBpIuOwlkkqDGHLOLAlz8RKq7ykNlUM6f2YiHyAVYhiRCLk4SPpcmeWQg/I9pVqt3Dbe3aShGIhROQmRdor2KkOH7LsOXL3LnA5ajkeHZg8deh8+f8hxP6N01ka+JPd0KGcq53dkkMlnSWeo/HlYd9mEPjff3SGZuzl/yivlscGWCgHVu6RCkXYjO04ObUx/MThj99oD2rS5yD99h8rrY9WtOBHwZ8yRtmrDGdHZSbvmvpf92h6arHXScyJtuA0ptOxOtsbjnzYvu6URRvD1sqdmK7T8z5TPMt5bEj+7ZPVkBuDJQtMYEo4rHbGWEMMIQ3sa9sQINugZvFrTuy+YWkzqEQyOdmZOZu4d0xQDS6SOm7w22tQ6nuVLzx6JOJtjzVj5r+eze99xrJ6Iu1jIEvcIngHlND2rL+hG7iTQkyNKcMtwBUDNiQyy08FLnzP37WAOxXkJfDY6Dc3RFOfSO6esM79fCI2VGhk3MQVAzfM9ZODetzGAJ3mkItX2qghQ/r9wXyQY017HzWoRVthZTMIt/p5Swrmcm3HA0VBR4Lbk3ozkZEY+/pz7UDUy0B4bU6cNP19wekFb8ZpGF28w5zPAAPEpSl2AQMDFsyGnvUWKVpfuyNUZU4eFE6fiJvlBbAa1mrc4DwDykiiuRUkMdA4mqCFQe9PZ4ChWSAN4VYKvIgIGm0ae0+5V7h2FgzGVvMhU9e3ULeqBoGLNwja6bI27OWv8GJiHihjSBCFFdehMaUPyFUs5JrIqNp5kErBPrnSH2264R5MlGxqivj8JsCGfDhJi4cHzRC85T5MwNiAy0YEmVIlAtFrYjD4Ao3bQvDLcKWXjqqRIFLWijkCKzF0ucN7IZUEYJcw23QMR97AGgco1buIZxqsdI4L1XGPlg5Yl6iLjTPvJA7GFYLYh1mCyFRbfQLMts8zWd8wIpiy/1q8S8NT3C6oLqfAgoIxWnI00FvpZ3T4X318XN1GeGJfpNF2mozJ+zyfyrpvi6XSU0gxoIJ5H8msphel0fMl1UqRHlrcF6TXQaKJ9FMSvSoRl8MPoPHnguobh0gYX3v2akV6plZcoK9NK45R19be0oXKWHIPQm+2lsDoDhlhbDDbePSpFsHAiGsOnFoTet3FjgTVoUl0DuY44U95G+D2WxWpzAZXOyoxs+Huq/XOj5DxQC5IvBIMG2ySkHUpLWqyEd0otclGQ3jVLRHszN8rIJXRtmGI2ouuoAVmuhDpDByWcexoq4PXsA4TOtXLke8WvquVXTw0ggVj+O9cpvpeq0mx+0qcNKMlrzcb0AdxMaTXymQDUvaNjVMdnfCZyVGHdYxplYBno3jPpuff2v4xXHFFCWO90fNqTyplrWvqO+zhT8yBeoe39f32PA4MNxfspYKlUbGknsh05zmyHt6kOmJ6HDqQmofGl4flz8XdranfOx+QTNaVToz4n/1M2zBdK3mJMRYqr8XxuDYKq9FSp27y/VtyHvdRzWMc9ZTLa3ndh2FWVnVNCgbgKwEplyJupFLEXXu+W0t02RIxOJ83Dw40MryWdA1niHKFH1aRRKGSe3YxyFrE96rYM1lmlHYOREKXHU5Qz6Q6Qw2oVsYJl9pifmM9MXb7SGxqgIqWUlKrmQIcZ0elpjax8q3JwOUgaEzejp9zYAG8JKWFDVFDuHMkYg7S6aTsRU1UIRNB1Z8dm67XmHjlm9w0VlB6dh6ml4DHgXul7u6lPQLeKLxWds/egDypbJDrsvapIy+64lKQ2wfmMUcb0XNvGRjsZtyozqhRkuqIA4+FWI93UAfeo4tmGz6GZoTp0sSad5djUJYDry8uucvYk/UOnAjjQD5EukYnSxxD/VVPY0tfhGE2p2FxNdDD+s8Ns2ROCuaoUcrAZoCdo1GB0nCr4Llm1NCI/ITiVpfVLa5p2pAu23Rk8tmW3roqT19+Hw1iIgDtm9+5Jaih6o7ooJVaS902xUDugsTnUjQkzirWWGLTKgb5mK3Ssg0GWd6RBChko6weAEKJw4eVYMKCL7AwcJyd1eOOBp4w8hGILXI1q3gHm44okFZUCLSx+jNlYpjKkI5QEN+6FGDdYn6WFXtCwovMBWOeELiMqLke3fMvwqf9nCA9BV0VTVVTkWNwi9Vp0JUN2UtoQjSNtUz6uQxt/osgnnkWk8nBdnmlQciEvkWSwhuZDHwgPerMV5dheQ2eH+n3L2r86eZGoT1B9TA3DYMPZSkOQTYvZFoCI8mo9J5lnbUJLu1IUZVqCgOFoI1JjeoSYkQE1tmHUANV0NT2XwTDZYR506NCSC4E7A6SeUXwRWJoVEmOEd0dHONxMg5j+iifKvXRPO4WFk1qoAK1J7OIfhbhBp4E856omBoqIy5sa1P0MuHef4W4q/cULKI/ygopdA0aZH+qKPwj6SAzT+XPsofBoUW5ZWpXc2+s7Oo0cEoHskmFf+poL1OsSmlT4KU9jemCCuM4DEwaSbLgaefSeyhv7MDZ9z+Di+ZpgGhvagjhsebDjsEubIt0ID5aIPr0bSVXPlIkOQbJgi/KnHECUNrfx+bwjNPkLPRMdXdzqNVR3Eo0EuTW1E2Vc8aX8q3RaA2kpQ84pTGCk8x28aa04qg0YopkT7ZSUvuTNXO9BAt+dk92hNZHkWAiI/Jn4i4biOOC5xnIY7nEB1IjKsh+C9pzrZx4ICEIcjkB+20QQ6FvApkG7gP31gw6y0OQ0rKPeZ5t2N8oH5FSCY/C0R5AwroM+15+ZHLrSiDiv3lXuXUqKkIGFtu8C0bSdYeaG+LHsmQIRKhiY+fkzvBs8FF8avptKvSESxqZtUUys7aUc9XccEv7ENOZYWO87LFCObmmEMuaRvImR+myoaUYhywz3YXqUNfS+1qOk8ZRqLwyuWGSkt+/YDAcW8KwkaIqzSKxwZHJWibKYInVoMnblfPq5qPZownMYTOhE2FiU2o8WsZ6OphtI2E7wFogp75yFSL2oGpXCkySaVzoiWW883w6ObcJX77vY46EyUeIdpV4NY3OSRgb2NFMUIdri+bsvvFIhHHDvG0ztkBOmnOdXOfQEydPN6jLgvEBIeo89ErC6IPWOfTy0vpBMpFmYhHg8yG0aVL2x/71v8kZ0pQd6L4chRs0tmKjzkUO2fP/GtHeHDl4ixJ117Crdzc+dqDpt+XtIolVObcGy0D7zcqKGAM1Kz5e9gdeyQPOa6GW8DDobHnvZedglxXHNoWqi0UHB4l1t2QmV2Oxwjw2ZkhgyLLnBSZIRFjuEJjyJHXX5QdCScHIi86/4W2SlGtAKZey1XSOMSpC0yBjlcyyb5YH3MirBMojoUm4n2BjPr+fpGVWBvPsyjbT4ByEuAzL65YyBrJLMe05AAptyhhG588ArhUoHjEA3hPU6EPB4Z8lze9+m8RqEYoIjACsDGmCkvQA0Y2EHR0dDlcgTWabKr+ZwVJk7Usea2G2YKMiL55vjW9wpT5/hgvsAx1jUHiciojOqZrJI4cb+HjnGOFBVreoiNFEXcQuxFbHL8r7Vs+nn1NIuQg9jMLNhzoiNz82nT8KdFyaz8pVzaOF0bjrMSsVk62WznrYk5adjUnokpOA8dyh71UCmsLGlBkd3Im25kPC6PKK891c9Mypv598x2pgPNrfAAJuzj0ARIyOlvPvQQAaPBR3JJ1UIuBhZUciDWuxqQnbHcEiUGrQhqldDWLMVI7gTsqk9V6XDKEtp4yI/5s1okCArRqHvHVqhhjR2NVSFZevwCMWErVkZGNHU0uPgwQTnxGov9e/ZTSm4LDnxBDH0YrCR/S+xRtK9ZKqlCg5awu1itTtTjsNcvyD4CkXo8Fs6BAy5tgwy9qSLy0LDlAQqkSMjkwGYKEPXn42qyTjecs5KZ4YOSX6vHGREQpHIvDS5y1k2uLd0gu5A84bWWlhj8jVEozZDVz/ogOc0b1dUzqQggwoQfFfXbWsAn2NXjoLfJ4cEWAbKMcAJMRiMpWsh70iZTc6Y6QI8RFPZ/6G1sWGfEY53bFGI9xm7d+kkYHSQMTndzai2bQwa/CwzygYk0AonqmBqmPrsPkhNMw8GqhV5QdO9jqNxuTzphD3HwdIVrEaDjaVOIQKXYbqgojxo5a7eF+r7O+pyYyiwZQ9AVnEQOaKU9QGvN7BJRh/VlykjSLxj922+R2n3xYpjL9JnjduLbQ6CM6JROq0ihrimKrkRpjLKN/O6nZsbPPYwZKMVwP4MXWpUU6CAjnFC0245JrFWWoMkFglzazR/GKdSnD7k+Fpn8DkiAopYy8eKUYbidnI/qSmRo0uqsee7ZJChAcfptyHVLGm8BgllqZR8SSA9RW1D3urGA6pUZhyxX0SylSPJn9Uf6ecJ0fvYjAege9mD7M5CDZnBMIwk1ss0bnFfKCekWaQumYi+4XOvYuYHZvRGp9938XlmJEjjvZZlncFlTAEDQe9Sc+G+AG0qnY6QepKhRUbozALAPCKKprF6hOvpPdO7DTV/fmizGQu5i4BvQTDp7wdcPcAObFIzQ+MLqrwVYiQRT/HgE0VZ8Tk9lzEjKv8sDG2Xf66Lh5pIS3Oy6HUHSXhw8TFTwcy9jtdi+eUMK39nVyWZZxlHGINGy4tQY28KJ4Gb6a7RihQBqZ33kXQag0MIyNqcb4/0/HR52TPg6ZxS+t1WdISrTBMCMdjA7jvXcmIZL9KnOC/6f2lAxrtBBVHzeGHS9+aMDrLziaIANSSmJ3K9SxCiCbtNJOhSVRk0gJPOPasme5+WwSoRYG9wVWus8dAGwRm1AXE7VY6sX0W9hrMV0c9nsENkaLUVcn6JSUJviGsrFWTnspUBzcUdwFQUw7Ia6FyPBl4EhGkIHukq40yY0B+7ehOpWZyvLhLVmCr5YCuZ3PGZVBBQgDQA3eYY+HKMgG6CJ/KaLG/aFISKVHJm6YV2ZO47mWv96timR4o7CVSz3+VngDl/9y0mDjiRF4yfW9NgItrHsyQtioR2PCQTG4IAscJI4kpRRVB0jyfITZ6AnIQ8CJeS9AMk9kodgn43UY+4loL0SkEiyo4DUgKiqK9BNftAPIq6LfPZ/EVeQtWqhIugDqHvCHQM5sCuH2GW1gGGhcTwCGOVWkTgCGeoakGUjMnOA4CpS3lhtJ8SZU3tgPtHI8YGQMeSVQ9xC4VmpB2A+2fNtox3kk4jHARdNRZfx7q3E1h4P4vSD+e6dldpGWwuVOWmyNJmSLIe1CvEd1dqXB244VClQpZTVDo88cqIDknzdS6cDgxQ9VBIRVcFKE0DqnsaNscIxymkCHA1BPoeQglr0ZGvVB3ug16KRYl08kp9yfUNRH1yiWjZWTxP0wF0+/UIk7o75naY8MXQ0JtGr08JaceSZEq4sxQZEK21GTsQoqmjFQOL6ysaCkk3piTOpi3NIZjaiXIUTFfa8Nz6FeQfy7QWRjrZKjYQ4hhISCaBGYulS42QlQJ5b5GTBLfekcTuWJJ0Z0mQ5KPec4CjgezV8q20pRjxPLRgLdycvn+i8RfRpea1hlIBwhT9GhZfMBnnNdKBTe1EoC2TBFg/K4K4cb3nDBhB5MW/x7iAKQ0qpO26zXxi+bKqHuV0RVoOBwXBvjcOClKpHExDBNOzzDgQiCZUYhNsOkQXshFhjY4JK6j/JFDqKt+nu8r/M6yLX0I6mGYTmni1HJUQDmJii78i85KkvRAtEoGmpJoIWMR/17oyUAVHtaLAi/uCBjR1Ea+in801wUyE/YSlH0Op1+h0cno6g4CuOpxMTjnQfVY/0pFyOpeCLhbM3Rc0X6BqB5LEEYES4qIFmvRd9e0auzXlBsev/UExvSu/tMyt01BQAiLNqYi5iMZ5A1bwjLBeteAqq1k+U+aqrH/XM1WU0s+IvNnXGciD8W3pQIrV1kAbMF9U05XltyD/bSQrxXWoaUwJ4JQzEyAEQQeh1ExKRI2VzxZo7wOCAeS0RsnwZ9Xc9Xw2UYUezzPJ6VsDukg4qz3K0u0mIneXBsJjtgZaHrLKwQ2wAcVZBRU58UgzAHEbC1SG13i4GMhkxgCIZW8v4ACaFKe7FC4VGViqxnLilp8LItvYa1XUkMCva2L4aK/iq9wHRJJmhlQ4D2SmglGkGUsGhkC/1N/wKgU4ag5pyhHieYwBJFvpVSiQKFCBncOENRPU6WxzWpqedxCFiSCWTUVgbXDEPSlzTEKeIXInW4xZWpqy/dmRXZfe6+/CagAKj4mOje64aO2Ahl0Hr8piUeutJpoilJDlnmKlo6OzpnOPzU+CuMtyjPLunulTEoJWx7lEQDrcXRlSPNNwyFRZCmRTqKGZyMiCckloJiOuGQZDpHaqELM058VpYB4Ofw1wCWPbwVq0GMdrhEOoOaVq148DGKVWwlsNpO2lZITv4oCREC4nR8LVq3KkCClyWnyXZppYKx1NrI0ialXL0mlTlWl8JzU+xU5IZUnCPA9wTzsJNMpxAQjuKZKEOdOWODgxDTsOBWlWpnGBtNgQCFajiG7dlPqUY9EeVYMYCeMBSYUDqLRcd9mG/SM/T0S+Bv1G5YrDc8eKZJKSyD3eI0sRaKPZARIdcg9L9iCkS8LZwh4xrEnJ0HvubZbl4Zh73wLLJg02bz0S4TYepEQVLRhwq3wyuhq3e8SKlG+TLwGtUGSkDocWrjWg77bppLqHiKh1CzZYLdBmiX5GWDiGA6VUsYhbOCGunlXSbRsdiv5+71h8nYcjFX88FDKaKENSabqsc1MxcXYiN8Gx0PCQ6wJE1UUDhPYOpyTqUOlzjKIBFefpMH9+7I6sC262WGzB3E4k3G2+w0L+JvbpoCIggCYS2UqU1Ad0qHtY3YIU7s7KUTp58VNGGG3pnNQZ2xKByqQI0Um2Rkpb651yZ5qfoVHVO0x6Rw8+zZ2duyvsqCUh7Ih32m0+CwGn+rFvUmCVZU0SuPqOSNdQCHbZIHomKuWQmCmca1UY4st4W1g7wfPoGUQWvbt7OG7uvxZKHBS6/k7Y67Jscp0NDcuyoZKXvFVDvJ+prF5zOiScUwBf1EWbvSvIdep0VLOhuaVHUbPWhJCWVvkoD2oeFENSE4RbsyCQeA6hE5JeZlOULS0UgcG8B7nT0GJ2hS/o6GlYZhMmO0wH4AAktd2T13oJbepZjbkmF9QkJpuhFt5Y6GKYxTVkGqEoqNIh41j4gv3SZmzsspevpuf2dLfp1pDfSkdmQivDn6YPZEQDSERrKG5Pg4kDOXN+R00wU4ViakCOXRly5dEBxncoEimNQRqhKhPNGntAmNLkHhTJ5+4krpGfrcOlVAOcPZHzUqQtIZqJHaFugUS7NDGOmKsZWhwFEKtbxax4FR1M8RJFPnquRZ4D6/lZ01BZEYII7oOaD3IGQmSx/tVIOQayNk1QRSNl1QjxIrgDgRbVSRrnSsN2ZU1hy8O9HtJ92GCbKI1Q/VQgkOR1uDaJ9mhvMYNmv3TvvWOW6aqhJRVp2Q3aMr+uGRQ0LZcGoYRNBTe5QCaYOKNhhcXXJOU0c0Kdejq4lIlY6AIapuwYHUe7KS+Nx48n0ng99XfIyJpKfqgSkaCrWcOiPNwjgjQ7oJBFaURFpCiRTYywnBvABW82B7nqC4+a5zup2jDJUfFISgSTDUtYodBRONqM8pAyUSRZR5SpD5LlFhoK0doKztECEpDlz+cowuKMYu9mdATxN6GQZU5T4kwEuOf6me4StZY9PIBhbgcZlTuWJCTTSfKwOT8LqbochHpQ82Kgr9hLoh/CbKVcI3fQoNQ60KBIv2wJgMGzJyfeFnm4GoOqlK2xT6N9wmXnC0uy7Fx1oUedG01y061gnsgo14GktsjGwFfjaEbjfs604ZY2Du0ttRixjjMWOmqzNiDQVdb0JjvA4htMdoCQoG/zVISDCqLZmSov1nzWGK+qLFAf4FERTwLP6ual6Di0fME4RC3LVsgNCfFM2NIO3sNRuLT3rrbo6NTUdYnNo2zqfUG3NdRQo7mFqc+3FZZ+DE3Q9mUTB2DQEARXGf9ckmAKkEww3NHVR0Ch1zLAcVUSYEDnhUDxfFVuUxnKYWmQMiqHLr5ByILJ5bizUck09BccXrsFWGrW8F1xDUId3jdkzjdMq0TwRhqSGarvwtG4QUNV3HdYMr0pxxTIiYNc3UvIA0JX72gtoHszTSPX8BoelDYxOm2wsDciysWcWcq28Iym7Iot4ltBR9yBCO7hYLljYgcqvEdnLYJInyYOQE5eQDxDCblqiG/P7wBTB6WvJkLQd1GdsxriPCKBeHV1EAdKFXHefce0ZIfsvZBToT2qJF1tB5HyddONdmxuM6Aj0ufetxzkFOuyLLuUCHRjg576f+h8u+9yji1gWMiD7OTkszq1YyC3JElDMLfYrMNai6foIemxZTmxIoGgYEUlEV0RuKoiId1/wGbV6oU6ajJU5EkB2TqCbFmAirjZRs2IxWeY7GCAWmwAtpkSYJFKoXZrPMRTO4zDCAN0kbExorYVJubzer/4ezJAZOlrYmkZg0Q7IkutjW7PEjMvzkJirMZ3X1xa/BDXxA9N0eGt1MAaRVZaS11jN+fnAoZuCz9nBbcJTZPKTLIsIZmafSC1ZaTTIQSLqkg0zsVaM+JYRK1dL5lzCPMkuDKExN7S2aSNWItyJiwd6rgmud4QQapqQkRdzZ8YpdpqhFO6lzZJ+9WB0b6pLwe0lXgWgwjYSq2AQiUtAhr083THpnb+4sumdHZKd8g/Mb1Gfl68a8eOqWHLoK0rPcefSXK5GR0W+TxMsFbnKRwauSww/+0g8ubcEIRob+mbKuUqy2CQq/trAp3PYTjMMVFVhzr8rV46pbaV48gAMmcaciEdktjEkbRaykElwpBAiBtG4k6/pJuIZ9llWpD5rAyMELnIObHfGr2nf5aKTbXwkNfGog0lNnjCYtEHS98wWtf9FKoUdL0S0QAAIABJREFUqFqUzkEkHXkHRQehm3geIoMYiap4EFGqb6OpCAgkwopUz6dBGjggfsRzsreDw1L4rrp6IMRpJZBbONuy00l6zsmwREtZiuTf0p9nRco9IimdDnIN81jnnogoBGpASzjlahhEOhTkJ4wXMtUTtORqyiGH7WmKu41OR6XmREM2IJqqDGTOLvserNoMA8IVB1dITlf/lWOqM6E9C5Q+DUicHJurS3WbDiIb+lxjA/b7T6ILuj4bCJlkrbNXaRsdcWWhxJhh7+F4qHJFLwSGsLlZhm6ogatmJNEaG4ToaWtCz5TaCR81EKZWZ+VgdBbDJGup9kTqqYtS92WmvWs0OZ1U3ECliBscS8LkzsM4aC+EhPTvTVJZwlrVnZUOqT5ffQQlHkoFp/e8kNYhQVPk/rrDspp+DD0dR3hmN3ZZMgBO0Cg7KyGaypEIhNfsAFlyhqTuI3cDpLQdanmmw1C5EyLWAnstLjUuD6WzP8SrhyL9G8vE6k5M/oA/p/RHhu3uxX95QPGqrtSsknDAvAN04aAXcSq5P0oLIjSaNVYO2LXZPQcedZYUxU8J2dIL0PCL3c8LnuBpa+hSWgoRkuGizXRVIrpSFsH8JfkfKW7NQ59QU9dYJUuHHbtRa800QOMIvCp+oJ4nUBDPj2gAl7XE2QlCuaP7WAAAGlbJc3T+vY5wctN0wH2TKzOia6cviHeb+7IzGy5/iZozIy7zIs+IuEDDYCXgCaVoWhYdxZJet2Ob1ZCeuZ1xclB5Wnl5rn4iAEGnuIu0JnKrryP+zpwVAjUgqUzofYlUQ+jGaAyplYj3lny3hEBMOxxQ63dO5MLCnFDOCAG51cnpVXDWS8kpO59VzVO2cHBNl1fXZ3bU9OhBzAYiqybUtgAiNo33WOTUbYmRdIN9HIwoqzHttJLY73cCl/IvSq9stzdACteeSkMQze0yEqqtXRDXSUQv2cfTsPDGObM5xtQBKesX55BkJKNIToqC5+yKCArxnQsqqOxpJCw4jdrvoaeo8RZ2WDr6xUvyL5GTNDBIcruG/EgwBjortRSMJdE4IFOUOEm2ZuQm36VJbuGMOAGfwbxEYx26lCqC2JSBc/EtkapzToUc4AK0lqin835cIEr/pZ2SnVAUl6IvYG42u0pRMLVMOzS9CgiYFoeQRJQ5ciR/5qohCVUjlw6KxFa6JyFH8MV27+eVEBHl6VRy4rKY+4HwyrIOo4/ku1qESnVIaHJB6xirHV8bVQrHMSfO8lvW5704G3I4WZnAOAk7Nr8iRx/emSXajFCE3GTh9fMF6ZUGCEVZIrnum4x0+YSMzDp40knwFOU/iztIPQU+UzAXCYeEWOodAsR7qFStPRcaWyUpm3+vau3pJPReOQcTtCsAeTUfQnQWqmEM3E6v/B7qdJ0xlidVmYiTQAbCy3ZqkrrtIcpJ1YAsb2pyVY0I2CNik6QeyKu9yC8R1KDdMeTnjz9XaYsClvanI4f35KUi+oxC4TDW2gZnVaXaMQ2XBUxpxzo7msJuSKRns3s35SYBz8pwRfv05CAsX9qg5hkaXTvgPRfOBeGf1P/EojI3jIMVRNhCSJ8OAsohVWkQdclNVonLUZuVRiEVZJS0gnhj16W1fBLdGxH1+Wqs6fTcMmopG4WywFLg4pqEhYSzcEebagCODmshAEYFObN0KkikhFzvgQwDEg1FIDO0IWUJ5Z5ayEtm3NBYiRpUqlzjEUJnbwqcSGNKw9IcTI0I0N4gYTryvRRi43lZWkWoQkVQxjqRH6CT1eyK4ps4Ot9A5W+QyA2ajBGfGbxRlKm7qzVBkbTDyOSne/NoeCw9TnAzngR1pavjmhmfGYT/NKAMACrJphrVgdaq/TsJ3LH0n4h0ynWVzsK1vyJ1+Twi8zs0yStVM4wfpkfLABCoi3acp7KCRQQwNoNqcJNJ/yQh2wJvS7Soq4ttsmrGKi9qzGW4SR4tYSXhlQKxSqixNZzsDJVfe0L06nZrcI4t61azFzrLgqNwClA5ki3dUqv14X5JLbjpgCldiBQq1Xdyht6q7KU27BSq7Gqj3ROKZcMaD6Tq/VOrCkqKv2AILgPp3KRLSP5HPojrUlUpwWg1jvFwU0bcWs2GjKa4SkUAltcaDxEVgeIg4t1q4pUINj1fmpNLFsw7VH0HtINCQiI9vUhKHdREfVBzUvx5ODCW54e0TUY+NoplOdLU+k7C0sFb6aOECh6auL7PkBoH12cqoASSgIhLcTsVovadGQCITLeeCDKpZDlYgJcPgTNKndB+R1S2lFMwoARqNcfC+b7dkAi5EEvJvUVGWpMgK1DbwoNdfUxElSZ+UGa7QIJJcYgGdrZSlyFHWZd6NzSbnBYjwqrUjxrioS0Oz6NmMhJySW5G3hy/F5BRcyQZbGBumBCdnw0rGswSUT+nRYnIm9M4JE7J4SVgZGU/SzwneeFGPkAwFFHpkbeOc9/TuUDiHx5gh0XkNf3zvtAnDLpgpbo9O5Ya9NNZaoPKa3KWikSAbrAOdFOTyuIBDSIRg3SqLtTkB+ik6RYg7UEI2ESA6mjG308kwhLgCLkVoaD0Jv+Xc0Mo9hH8jqVs0LEJUVh1LCa0hd6f/957pqFR+WmYGNXHuzudRjwqVCtf93RE1c/EdDh/L/5Os0NIP6F0SDfJFQ/CeSt9rR3gs7MxToR4D3J8spmrNeU1FU32q33yjFbcBZZnM9VRShnfVr1VEhCGXXc6tOiSNjRXetf5npbIptmK4TyIcL1JnRkhEInKuFcMjg2asyKtB1HjIEuYe9+a8bbylMhSsjwqAh3D5ccZUYt4mtCi9NLDgNWkYt7Qjb+XJZpoFRdjLoZYTH5AR3IQJBY1qhxQOVPai+IHRD5GaVct10joXvmYcjrLPVVqpEWdKHiqo6M/14GoDVAvgOTy6Xz1yzsMhdrq75CJpzEbp5JHu3n4caVo8TlOjmjGkFCh4GVVOzKFU+QaDlseuuFQyjll6XEoI2JYu0Jwu4qYiKasDg8iFEA2TjF96b4LBl4lWQPct+gIeK1n8UXTp5SOIO2uxhHW5LIlvgq7fgy5Tq3VYmva3Y5/NryDRFMAdpyFgT3F47AebgA1C07tSXeVzAPZyZ41TkHDlOW8svIx8G1VKRMyrtSwp8NjVcLr3EnPNKZ1cU5mbpmU1IYxcGaA4ZlSp7k4FF1ToPOx31Ht1gTx5MFl5qaXTLKxZN+JQNJUWVocfPP+5cHSYajXZMh9+atBJGh5wMZZBDLYEQHpuRJfQZyKcu6qUsjgdOiUSysS2fi5NPI9plrQPYgDqEqiQ5CXAHnPz9GzxdqFbDqcqLgLvZMkzOMagt+nZyIchYRLQTCnQaIQyajnT0LUZcQYfhF6O7IpbSRRq4QLOrsqne6VxVFVl7IJ/ZsQXE+MY7QDVa1UMgS8fnqIhtq72qfBQeda989CnmkxjmEfpJf4DBtWeggbnqVV+mNTogPkHoD70vbWuy6rluRevUkt9xD5/UjILxQypspV+o9P/+w0tw3vqmcHsuKogCxHJXtN+1NqNQ61Kk2IrrZgyubz/uKyUuHbjFNKA7RptVBldPmyaah8MObBJSPXLIdWUmpoLsPC/HqQaSs/pCftkOJPuocgwCR9LXEUy1pJcMb77ah2W2xNI6HsFj0Htqiqkc+A/UO3YMuDp9JV8RtxrpaqCmX1RHd/sGoDjaOXQpGcDjwnf+VmO8U2w6aOBGQe1jQUTvpqMUpQKDGkyjuZQSABHzQLLjP2ei9qS2CcZQqmJvCItNmUpH6XWjWhVBFs+axw1O3ilsYvfU6jzqJmjZTqlWxtOtU65MURNVc6pcnjg1NS8IPn/pSew5jfq38kAken3JuRhevMJjePVGVqJ3LfOgaBmy+1nsOzLL7GpMFLJl6pFMNKS9wXTDhIDUvY+zb23g7SfrWyoQSN91pcVxuwOmiDE+ksiQ4XO+v8qToXvSZGFBW2NiNhv5RiLSFseiR5Wsfw4QR8LJtqIY0bFcBL7oSe1BklUJr/uJO5GqWqgWsGfA3BqXA6+xJcgaV4Hk8Fop4xPXx+5lTvx0fuhPljx2rm2Xr3QGH5MzGubkBWxoYr77DGzloXjJxDIOOMSUzz9H3JWqNKXemA9X1gmpRl5SHJ556IsJKSMT5xgqNul6+0qQ8gTXJlobHx+6NpqQhu5OfkQQOgQTVAzUQQ56NuUtlHEqV6PyiSy4o8ZOaQWK5UvjBAEvlIe3b5HSKga9ixBuEoDVNK5umEhHqQSLeqBkpPhUaVpsWzMBlWukvkJH2MRHBKLaOkG810AMh72CAzUFB0pheWwj2h7AH/IjptRdQLZS75uQo1lbbTjsxy1WPNOXtUZ2kwOxH28Gh+XNwxN0w+2wo5KQskTfjybXAcXZEBlWZoIbUQYIRq+bgFufQaigIFJcNZLXnXaix6/HcoHw53bqq0m63u6FnilXx8EQeiRfMdujc0KwERnOPo2QPhvuPFNch3FcpRRPIu0VG8/ziAZywnR46q4T41Wl33dUpJaGLaEV2nOe4NUXJ17nZ4eDLdWA0/g5wHodSkOyj5pvzYIr3KS3kU/aGRasMN5VaHu+T7csI8NFZpTMJ9kpUjIokgs+ThqEFGIudoyPl7hV5VkYi/oqobm9JYXZraDI1JDIuL75gQLQxjEKimOK3bBKeQraeTkZVXwBkYJhitLd5TgUxcmY4AK4VaC62loD8CHcYP7IsAo2k3W8A4Z3RBN6YnQ9RP9G2aUtbRPByAe087pvVAaY6eAeQhOy/DGknqELXSwRqA1m12dBOhyG4pVI037T4Mxjmbom+IIIqsKQ9cJTrBLkApiPJLwXoLI+Q4r4lwcYFSlOrZj/H3hSAKPUh/0YbfNziRyyIZbm3z4OxaRr5YfAluquYtHqA4DlkOl9VseGcNOC21pRBFOsnMg8emq/HZKNnlJy5d0mRWXsQtsRNYMN3IDcVezPndkZIFZ5E3YemAQ5UbAEy1cmYj90hS7+IWGmxAC3qPcd5ClEeH9JQ75HTMedFP2tw+vyT00dBS8SnBW7gEStCZg8ceqTQ+7+1FNnxxdd13RFw2vN/AX9jY/q3O0cZXWdKxiBSGOzlMVagaYHHjeefkWR/WQbZVaz5wQ5kumbJaAKB0W5SA9q00RYD0FqpAVbt/pl9pa8XbJMoH4C5tx4BNXIKxSNVm98VCPJLmzcMpMxqHuCAnXi1dvQCKGjKIkqHm9W5AwT45Di6gW0RmecuOXf5ctMSzLTcbsBrUKly1YkIsV2/IuBjx3fs3jw0t5HtxBPx5dRqWipGWlIuoJqBx5N//39a5JEmS5EZUYe6Z1XfgQckr8KLDHTekSE9lhBu4gD7AooY1MlJdmfExtw+gUChghWJOQzGIixnEaJLd+cij65R154xXCK3OBR8D3DF9wa9+7anArLmKlgJfmi7aZ7HWcA670dd0dVe1iMzJWKANUA6jNAVMdiY575ekNxL9rDL9e/2l5/lbVFpu8wpvh6GyMXgzlzZk6e9/8kdVdv/SiaXfx328tV7el/aszPu1flWflfjy+OcA032rJe56dcsA1onyg+IAhsyGN5OkaWFnBBHnvOsPo8pN8dPvFa3MXGA8xWfqscJtWClMWO/UPWrr/BhzoXeb/j5PTaYq9OxHO5+8lZFnnt7GUqS9lNk7vTeSD8Ine14LR4fu1kAIFuBMK8bAVoVWuEOQvwjm/DwYVLrWAaucdQxj4bMyWoJOg8KNcDt4YFmHt2gLDQTOFO39SE11H0iPa+nSHd+lxe9waubjRCfPIfDCYE4uns1PsDTZiI/xybl+r8CK8ZoYxhQwvGpqlKzTFNSdCKned2osPvctisT+Jc1rPp4lLM9+HaKq/z9bxpwvkQq8tBMoPX01qyfGHxmRfk6cV4y3Rhcj0JsrPY3klkPo+j1x+yey4eYyhH+90p2xGS/9weHwHGKdrjKXOB1/X33XPj4HTkn+zdbZsQ2kezo/0DbnsGuRjlAO/Ua4vmQuGco2eMN+SFf8UqXbS2Vrz6v82MvdqXengGqxqySNRYLAOjgG3jwWn3ROvavz8OmsQErkxQeKUd47cS/scxuuCD2HJZ7r7ioVyS1inx2k0hNw6X3eWJ6fJwGOZWBXHJtTB5QtX1t7cDe0q81ntJKhSzSlXR1XyqHCzq2r+01EcwAZk8ot8ZWvFjwMI8a7K2aj0FaLkTRZofBBgCw742U2HIanJOzVgUv2cK13CcI6MhaTGqxYnHoNKzt1fdadGNpWx7JRu2ZuabGPhlimyCy7I9YnocphYD66EPtIU5ezANpLn82Aoo2QPuYD47r682jBWN95alveHXbsPgMn6jS283ecfMcEHqlp2Kv+/lYyJ81z4HiqmthRksqhjZFuYaHOUE+9d+SwhIRBC8N6PkkVb89CibkInaYo0zUtqbwDzUFXVk4nKi7PJe4iw95SWW+rWgDMhxv12iPXZiRqNxHTh1hq6EuaNErQFVTOOb3ThI6cQTg2QZX1YnnVaTjlbDb5eNGjI0SqCvRACOEshq5GF7VwXxpyig12bBq8aW9eFKlr5qJDn3pJcQgju547KNXrkHo6C8JcS3HMwR6jaCSHknOZ55FRn/y5rOn7qF3AICA2aoSj14RwHnOHQ3ghDrWItcmktblX34LVB3Q0EW1g2VHNYSyJdKZDscsGtZxkGdjraIlYHtWCu6Nj/Y7KItT4qVKFozEy7kAKohNP6znsOVZ7bAwtx3+6scWRmp4z0Aa7D/U87xkC1hgJ606dy6U4FcEa5yc7iM4SKZX68s8fLX036vrXzMhqERyfU/89yPLOfKJZcW8srNWp75+HuDzpvkEJllpAMKzUY0C37LUKfSwf4suWbmuXDXRPwPLUNmBJ497amNOX8ICnHVaQr6dTch2iS3T6ng1aUBIvT2wNEXZ4Bc/mGAFDychqHLPOfpR/QmONkcit6Tx26AbEv/uUNEnbXESjBTZWeh7DiMJrAPEp6e15q9AF/QL8EsRtTGVlzzP9MqO/j8MW4V6lNtKU5LPeA/PHMaTXv50HRh8eRYVcVkxasoV7OdmJau1msM4dqdRW6FV4gQzHoW+Rfz6vJZvkECsm40ez3kED9Xfpao7Sf6mfLbV1+2rBrbe4NmNkAC4VCM7E7tCDnTUhB6flkGv3PNMrxSGtDU47Fp+Vmhej5AMFP6oWA95BvF0IECu0dCB3SNXHGNXT3qldNsbwqmAYDDQPMgcIYU+JVT4vRi4xybe43bvIJ2nFo71/a+uAtCeBYtFI/Tkq/nIr6TuoA1FwgIH0MqGTo4XHq1Uvhy/pUKZV7Li19ToMyQHXjyeedeXSYCDehC7DBxR0fHL6dgzTTpMTCCDD5g7fjlDvMCgTO55GpcZMkZgWEFaD0HK8S30OxPHlOS9ScDIdeErI2+FckkOnrerP+BiBZHstCD8yOU8XEdJO/9GlX9rductMQj7KfaTRbWLqv2pM7/1PHxzD9VjuTQEpbCFfTgv9viM1q39HWVZKAQpuN/G9BlmdaWHmemdKMajhArHJcnyLDosk5Yb79zxTStwBvNushtDh8Dpa5hHeVcZoEFhJvU+F5W4BFw7mdFg1D5PKZ16qcPLLe5BzRqqX9PBy0uEiDoobn82Ayk4drcgPL9NxpnZ57CZCLnu7Sf1QR3FZRDOHpggxsh/Ayo7L/ZorvkVn5yd/uhW7hGUH6nKAjTYcj7FoRY7zDM8cdP+dER+fSygw4VFiPzpNSsPhgYazyU4dQSi6gQ8c0El+wj5XodZAX+LYppVmx4ny80ZwH8TrZEcmpRyNJCad5rF7/QiVZn0qtfz0PaFswjDpPT+tz7u0QD9JGEcql4up+d7bh40wEA84Ha7OUG3QzhS11XLsFi5dsUpX0uYU1HN25J5wob7P5GIM31B3+uYxruE0OBMp8BKhH2ihPDIhO2n54m0wrKF1PHsJ3movsg7KKe1fR/mFNFwZhpMaIviQ3ibMWyzv832ER2o0rCadWbfhP3DMoJnIyPsDOvtFEp4k2rM34TE7U50ODSkSsvGQInvQEDkggEqNlTF5ko7cE88pp+isoSuX3B6QTgl5Q/kv/IE5FSv7znLuWvAyQJfoKj1hSgikQKigttiDbHLy+334JeTc8zoMyuE5aumYwfYsiILksKUMmdrLSOnbyAm1ZkH3cfDOlCdh1tsXT+NtaQFPp6inN3z2s8ltBis0gIjc7Zl0HAq86Jbbz6v4lyLL3Bg4Ga8ldUZ89Xxcg0Dh4tnpag50W8UEl5wZN3UI1BySER8XBZ3ahKmpGfIWVELJAmtXhnX7QE2vFvp7ci1iobzvRoaVImXkNWeV9j/T4p9niZvQa78crQpdIkEatJDMq5+LHhdzT8kQuXxRF9IJlUkqj4vBcPJqfYX6zJSxsjWB8Dn/T5zOYcX6VHgBhB9+g2xFz0IyCZRCDzHavQza8px1/MTn0wGIhx6Vc33BeX8CsJi7FtpK5h7vamMEd8J3Q5g2aZqWDyfpxvHgU4i2hnA7NuukHMdKI+jpwroeoxcvef/hIT2G6lB1q7sfCVHOpLgwqufkgzIu0VWdw0GodfIL8/pOXWMk04I6mavxKMt41OYnTq+itCmOGgKQwwYyZO0R/22HRpNNYO9wkLqw6fg3lcmQi2eRH07qJBYxxpnVAwI90DznfAZIbsbCnqiQncuYxPrLWb4cHNX7v6tPD37s2P+z7jMfpPH73y3a+te9wv5hz/bf7CPpj3WlupnyB7u8PJmUU5eUcW8KnxIIdlwmFHeXoVcbdheXKLoUuVDHHDwumWlrnqc4aIgbLl7phW9jA4se/TmzWOlFYrNT6HMd//7RFb/83j36iJpxz+chskpJTdLWRghnPljUT3EZfExxHvPdhEVwK5qfzdMIQu3Rj197ciQHAjsO6t7T0Zm08mf/UngbDCQajDFWbGRINyDn6B/yA6UxonEQNtihIk3pOm1koYa1y3PsMm3zQ6l0al6GwfWa3s+N3upzOv7ubMX+IyTz317PESsVAVzOZ2T44b1JOCOli7kORxSjR+DagU+k6YPnczG3oM26dSjrv2notOJLNCSu16J34VnBdZTOr87UVAhPywG+C9Q38oUxUCNAnGV8lC0xV+9T9f5mn4TXDRRFaK+8I1YW/1AHnnb2FmJoYs6n9QL1NQMjZajYF9KKSlP1AuOde/Hi0sl/lJX7JTwk8W1vYsOrmYQwmZaaawhDEb8El3BxT4l5i77tS5NPfnwIV96ll1AdsjN2/tAzBO3q7obAsyIuHGsj4RuodFxr0GjLiOUo25eteSTp3aWt1zGWSzJyG6ER81pGoJjzugOTHDvrU+tXYeLV1w5sjeibMQGdsz0cdRXFk8jfCLfFNX9ymOixRWW93vrRcCzptbl7c7PmhLt005KmIzi6kGlnbzYmVmd1zh6r69BLExIybzWvsoFLXfFL7/xnPZM7m6XcHUzZ/Ne2E2O+ujGTbu2o6tTh+zxvZD8OLmm1XqJCoqIQnubE6jPopr96bko+ec/rAhJ0iU5wl5s9qcdY4i5YrtqA0XzGcFX+k48qXX33+cMx3a6/8YfWhkcEMrG347R0jYZhZl9hH1aq5aOrY9+Re7e1axITC41VnnhuDt/Wc8TrW3TePngDvUTFXRmgQSX1/Yf+QYNgLsfjO39ENaNUCKuhZm8vPIhPup+vUNZXPwMbrzqBXT1eQaBathsilUjRzmMuYnQZLXZy3B95suZ1gB/5MmaNwGhp9ffWes38Rl6Oa7dOfkCS62ein3kb4jaPcjQ+yjiMd3tEUqGgjombK+e/+9/RBnMa13bYoknTyc9DG/wzNIF/6dBhPVX2nuo1mzS51NAeLoNXeFyUl0uDwspo1zh3Sqvj3xlfe95GT2W+n75Cs7J5fQ2m9z2B+IlAcSCVuWPvPlJyl0tIMUrLUg9PBqlv69sv72F/skvhQXjScC0gyKnmxjBsAlMhm3j2D5eAQjAMFMHGYdEiKonDIi8gi5xyQbJNOCK5X8HceSFN3PS0hxwDgrdBYCPJxI6b5BoHsFkYId8Y9rx4NpAFJFsJz1AJbndsnoPO+8A1GJpmoRWa+zUnU0GKL5W6jK4ufanviNXqn2MwV3us0O1iLw5nja+29+U2a2XQh1Qcg2fYbN3IZ4Ofa46dS+PP7usfCtYY7IdXVQ4BO+MGIYF3Do8lbOcY2mlSOwhHPGPLj6egqjUfEOcqb4pW42zs3KRlHw6pie4cTQMirHJqbNsRSVXm5xFB0Mn9NI5oFTAIhXDNKMnSdZxbq4tzfcwPYRZ6ilAocvKA6CLC/0JwxuoUAToNosg8pX7qmeLcJ15DRe8BQs3P1Rv5Q1pXwu9r71c3sxtC52nWE08YdaUeU9gkluMZ4rG2xL46nsyDPdiTb20TYbiVs6GGdGQJnLaclmWUrj/K/N0HZeutt7MZJ0m0PE6Ya4rSJCDt4wn76fG2odRkKYb4m/BAPT8zDxN+mOeJuYuCEET9iY5No7IvcEP0PTg959TGyJuhMgyP7DVi6zly6c1ZJHLmyuiXYH7ax+MpUqkrj4pcsh3eILRu2/2ZBcsrXDNZ5tRq9/VozYs+ngeSbmt6eCirFmLp7uvzzv2Aw2BvgPj+hMyTVkU1/K77QFyysOPpMUGu06O0RgDKrXl/BOK7mr8gfd9ZNu+FUhq/Bb6AW6u7ZJ6a5aQgs/xRN6dROVfmj7mb7MojyNNtZNKhsE4kFt4X0y6y1h9ODkNczzcciz7OzaSht9GsFGcbByOge8UVxFk9KX/m43uRTHT6ot+6ZXusXoazDraGj+PNvqE8JpcO+ckdnGPdjA7ydm1IeeWPOhAtXfq2FTZ5elSA9k3eboyLbD3MOyxDs9WHf8jMxiktSTcf0rA7On2Zi8+eojVEamVgZe84SIG4djoZEcaoN8CgIAI6em/w2uEVii/46sNU/3tJuY6cPl6NLosfAAAILUlEQVRkei7UertBCygEQlh0iYbAlDBwo0RcosISJAD/wZ7xqVDqrZVXP29xJrQI+K5PjTGel/tTDAI6yfcJOZFTh2SysniU7CsUo+d/NZ8yfId8eKpTOOll3AQFW0isOawguKkIpmHvaSYv3Xr7efhz6etjH18N7EvE1orS1oeE90uK8ndK+0+NCjoYiNMmY/v3oBY0GXP1B/MLx9aNe9zF7Niaee/9xOMuxsBiHqbml0zGMNV4431YYmAZjTSUMkP93QsHfNwwsVHhwJO/TUxmq+3wCig6dyIKm9h2roZD8AS/grKtDsuT4+m2N+4Zt21a5Wlrt/p0hDl5zBgt9XY+0v5RBmrGUVqCLrybhJhNml4NiGvYcOOJ8e5u05aPOxXh2RjPwNopi6+fYYi2DWHfM5GpcFf1d1T4lApl/hZQOZNn8NzLoUMz5LufkVh6J7Uf0c9Ta383FwNBTMsB4PPOly599+1k2MwKX8wpbO4RieYDat2qUJEQcee7HBZwu3Uanjuc6TkmgV5eZUjQkBzh0M5H9/rlbf2H0lW1vvJ4rvj2mr97/VhT5pXMFRzVc/TkWLH0PsrQpwFQCuHZ09mnQXUjqVfLGujkXvzfqxoxeYXiGONZp1LnowjbDj/j0aOfda+4961vqSWuE6+vZuQrLnv0EsqzgUYQmKk7/ppNF6lL3+NBVB5Vcr441T+/9O1u2q+GqhfNWrQkq/bOQinQxOSvgcbFaFd95G2bexQxWecQlNDHZE46dagjTdcpve1NNgTp7cxL6FXHJmCyx8tI4RbulDlHHaL2SKs3fsW6X5r0bYrqWDY4h7H5HXvJ7j2hQ92npRVbjx1Bd4MK4leyH1OPslBDHk2LKpNU1OgdX0aMlw/zZ9YBIq8yYt+CyIUJIyWIhmTptoaYPRKaYjd3po7bY5+bwHa+mxda+qW0tAwtQpfwR+2wgdTshDkg9XR1yO/4/ngm1rPQTYn3Jk1J1qWUwFd+qipZ37JYy4QzPMwyzZK6o8ZfYf+lL38mjquzkjaCl768/sOxhF9PzVWNFcT16I7VNAOJBJANWiHC2Jasd7SxtPPO1eGFmV8lLceiyb+uJE0La5KLa0YlQMFW4PVyioUgvMLxKhWGmVs0b6X2YL7DcCxnMtiEII44hCkfsV6qYzDotPBGlFnz6iZeBNelq18BeojqTuI/2XN06arsBGNu0VaRYOFDIPQRftazZ+dkWmaeFsYUtj23pmw5jgzV4ye5ei6rEO/LBtDcQc/x3BmCGA1jGR8z45RwE38mtvvpGNP2Ky0QS2m5RT97pRKV1VdjSv9nH0x9Qwi+pYnKY/981gnNz3j/R/2L56fESdSfhN833w8fU++vFoesBXPH/sPjksHheeuzuK7CUL4zT597uEPtP/Zq9wTlPKQvTPJ76a5Pdog9wGvojggZWcHj3avV+/nkwHoPHNeJeswnVFCfSQRlNV/3s3905esos2VLPj2Fc2T2UUtRD4j12wH8cVchby46Xe9OIw5bPRLWd1l2qSenemruhu2Xi4L24XEeAV2HTCto6bAA4UzURLUXjqefYS5wtrFUFCSlGUs/+xQujUxZ2tYNDAF2tXdnE2a+DwAEmUW/B2cCgtSxBEQfHwiBiDAqNcVT1B3kgJlMddHSQWQVJC6icjvkom5jNs3q8TM3Z/s+7o8hr18TDyGZJsr97yb3KAMc0rc8JVhj6b1/i2if4qnnGD9peEhCZgZB0WNSHSNUz+imvn7asy/IGYbUPjjT4ylUjdOJbUhzuC/WLfer57DvrvUZOO/Xqacl5BzkuTWlENHSd4kQn2feMc4FvoYrEkcafiqm40CkzSJp6+27Wh4/rXvCalLYpM/Ln5rU3rn/8X19a+kqQYeFV0slUrriS7d7BuBR4ChG6lFkJ4VPECTqWBYLKH8OJehDJo33c7qwrdt4DjxhPUMcBVCQNDZovTBq73/G00cf095geO7zEEoTozdCkBfmaCbS35GIxrKN0Sk/lpC0n4eYg8dBGhkx7DQXJ/Xr/X2T/cB4YzDJuEw1bcFiDvtu2XkbGhCFDbXOw5Qzn3g8bimTDfAdXw27Q5eu+PYeodO1V/rYY9P0qEjGy2Tn8h65vCfZh+U9q6oVIR/fwfcvF6qxPy59ax2fMVL96NdTaHi54I/CP9Zh5gWkVWEcyLfvyCHTYSNc7z8qiIValiBGrXHgd9P3Yx/fC+fDxh1UhtNulasqCiAjCZo7DQFh64Q4GCocJgi43r+W9Hr//V/336///ve83v95//XXv5F/3XpCPYUgDg80lMpc5ZXuhA1+YelV8TyW/9HIodlcZWjT37GqM2Ks3PlExJU733Eahuq+OFLVpeJPVlyZ0lIWbbTiCqdHd+YODkNGZKbjijC/nNUw3wsRodVJtlTGpTszdkau2JGR+WTEFZK0MnLHEw5XcjtFWUzNnWPDvdiOPcgs7NghSe/83zw3Tg4+VcSK5LlUcaNnNEKR1/pScXYHmUoCR2PY0tjnAJkmBL/06J0hRdrjpjKWrtx6pIisOTT/EsrMHSuuzNyx407W1eRc9H/rCD1mDAoHShjgFXfufNapcNA51l430JZ7M9RcZGqvpSsfXXr0DvMSieK4uTdRRTwtDupIP2tp7RVX7nxiw5Gw5yPz3EeTY+g2UAU6YmVkRJWrL8/Ple98xaVbYNesCwyTAytVN44rvnLnO+r3kbX2jp96d8hrUFsmItJZveU9GNsBMg2vC/GvjFTsyNi5M2K5QffVHiByEcfprVcsXXmu+3v//Y+/X//zH/8HedwnOfc+BvUAAAAASUVORK5CYII="},{"background-color":"linear-gradient(to bottom, #f4f4f4 0%, #f4f4f4 100%)", "background-pattern":"" , "items": [ {"x": -214,"y": 97,"w": 878,"h": 212,"type":"text","text": "","text-data": "UGFnZSBUaXRsZQ==","font": "raleway","color": "#a10705","font-size": 28, "font-style":"regular", "justification": 0 }, {"x": 1534,"y": -153,"w": 253,"h": 392, "type": "color", "background_color": "linear-gradient(to bottom, #ed5353 0%, #a10705 100%)", "border-radius": 0 }, {"x": -209,"y": 333,"w": 1992,"h": 638,"type":"text","text": "","text-data": "TG9yZW0gaXBzdW0gZG9sb3Igc2l0IGFtZXQsIGNvbnNlY3RldHVyIGFkaXBpc2NpbmcgZWxpdCwgc2VkIGRvIGVpdXNtb2QgdGVtcG9yIGluY2lkaWR1bnQgdXQgbGFib3JlIGV0IGRvbG9yZSBtYWduYSBhbGlxdWEuIFV0IGVuaW0gYWQgbWluaW0gdmVuaWFtLCBxdWlzIG5vc3RydWQgZXhlcmNpdGF0aW9uIHVsbGFtY28gbGFib3JpcyBuaXNpIHV0IGFsaXF1aXAgZXggZWEgY29tbW9kbyBjb25zZXF1YXQgeg==","font": "open sans","color": "#666666","font-size": 16, "font-style":"light", "justification": 3 }], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAgAElEQVR4nOy9d5BlWV7f+bn3ee/Tu8rMSlfpKjNfZnZP9TQwg9GEtOyyCyyCFdpFAu0otAu7jCIIArQIGdagAAKBBCOMdtmACdgQwo4RYnq6p7rLpvfevpfueXvN2T9eVnWZrO6snnLZcz8RHVGd977j7rnfe+653/M70mc/+9nv6Ovr+2ehUKgBkDAwMPhAbKmUqf13fjvyvNKPX3sjfTQ8nH9e6T8lIpFI7ExOTv6sua+v75/90A/9UFSSDJ0wMDgPaizG9m/9u+eWfueVK97Rz3zG+9wyeEqEELWyLP+8ORQKNRhCYWBwfgSg6/rzS1+I55b2R0GSJAKBQIMZ49XDwOApEd9UYgEgSZJkftmFMDC4cAjQtG8usQAwxMLA4Cn5ZnsNuYchFgYGHwFd155f4oZYGBh8XPjmm7MAQywMDJ4eYbyGGBgYnIPnPmeBIRYGBh8bjJGFgYHBhyOMOQsDA4NzYoiFgYHBh1KZs3h+n04NsTAw+Bih68/vhjbEwsDg44IQhinrVUaoZcqpNA9+VZLMFsxeD7Isv9iyCIGWTaGV1CeeY3J7Ka7eIZWwU3dtELQy5UwRq8/DvVW+R1/5D0hN44Q6al5U0Q2eAc/f7v3ckv6GuDBiUV54my//rR/G0dZB5V4TqNksvmvfw9A//8dYrC9OMCQJ1n/pc2y/tQaAnk+TXY/h6blXNmj+if8LV/otdlZC1F0bRN38K77yY7/Ft//Z72O1Vk6K/eFvY/pUvSEWFxBjIdkrjq1xgE/82R9jswACRDnH3Of+ByZ+4XcY+Zn/nhcXl0Oi/af/Le0/DSAoTv4Vb//DX+GNv/hjLKZ7p0gg+qkSRgSAjx8CIQyxeMWRkGQZSa7cgJLDS+f/8lm++Lf/FeXP/TBWqyC3NE38rXco51X8I9eoem0Ik7ky6hBCUNpeYu8vv0w5pxP+tr+Bv9HN9p+9S8t/918hAUIpkrxznYPrt5HsAao+/Z342uofEyLpwVcfWapEBZFlpAf+nJl6h+Sxg5qBCMu/+Ueo+2ss/eL/SfDaZ6i71vtY7YTQKKzNE/tPf00ppxGIXiMyNojpvgIZvBI8b7v3K+rgfLEv+88ByWZHqApCFxz9yW8x/5t/hKO1l9BgN7u//nNM/qvfQxcCIQTpd/4/3vqvf4jMsYqzNsjmr/4TZn/586z+7h8hAFFKM/uTP8bcv/sTPL3DuKpszH7uR1n6wn/+SGqfnfgqW391E9nhJzRyBdkTIPSJa3iaq+ER8RFCEPt/fon3fvznkILNBPs6iH/hV7jxuf8DVX01O883K4LKa8jz+s8YWTxjhBCgK2z+xm8TeP1TWJ0mwt/994n8l+/fhOGRLr5y7b+l8Pe/F4cjz+Tn/gnt//L/5dKn+5GApu/7flZ+7sfYzFXOj//Br5JULvPav/lpTKejl5pvfYO3v+fvEHlthGDTRwuLKDv9BK92Ibu/Tmj8NaxnzK+U195j5vP/mfE//AM8ERcAVd/6KRZ+8odZ+oO36P7BN42QZq8QwjBlvdqU9+e4+cM/yOl9jJI4QHhaif76P0KWJPRihviX/4KT2RWQzdhq6zEpJ5QLRczx98jYrtD4yd73bzrZQu1/87dZ/srvAIK9P/9j/N/5U6Snpx7IVRDqDbL3pa8T/Hvf9ZxqJjj+6p9i7exD3Vshsff+kUD0KrN//B/o+oFP3n/9MnjZCDTDlPVqYw420/mPfwqL+XTOwmLH1dKC2WZGKDnmf+qzKHWf5NL3fB8mi0RpdwWtrFfeMXMZTF4PsumRuYf7kwwCLZ8n8faX0dcCD2fsv0Kwo/q51k0v5CmsLrH9h4/PT9R/x9hzzdvgKTGWqL/6yDYX3iu92CyPP2HV/WX23z3mzbf/HpZTQXA11WKzV/5tvTSMtPELZOJZ/HWe+79TDveofAWTCQ6PknS/Sd//+n33Rx9C19CKJUxO57OtzEMdQsI3MIb5S2m6f+af3v8MLERFwEwul/EK8gphhNW74JgC1dhdx2x/6RYt3z6EcrzL9m//KumijJIvItddovtHPs3tH/0fGfgXP4uvpYrM5Nss/Nrvg+QHoOlHf5LdH/wsqy1BWv7mm1DOsPd7/5qN9/J84jf/+f2vKh8Jsw3tMEZmZR2zXsZzpRvZbCG3NE9+tx7X+HdTXfUFJn7+V+j9iR/B7rGQfPcrTP7TX2Pw3/8h/tpnLFYGHxmTzUZwbPy5pW+veTV9NxdGLCSbE2dj/aMfEe4ju2sY+pVfYuZ//0V2flPB0XiJ2u/+frr1Ism7S1RdrqHxH/485qrPs/CzP4EmrPjHv5XOf/Rj3PipLwBgqe1i7Hd/jeVf+3Wu/96vIlkc+Me+ldFf/jvIHyAUss1VKdsjfzd5gzhCFSEy147S/u3tTP5P/wB3/+sM/Mv/jfof+CHu/tyvcHvmqwx9/jfo+aXPs/3v/y13/sHfRdfA0dJF/7/+TXyGULxS2KurefNP/+xlF+OFI33hC1/Y/8xnPvNqStkzRAidUvwQW3XVfc+EEILEX/4Gd353iU/9/i8aQ30DgyfwxS9+MX7hfRbnRi0w+7kfYeHzXyAXO0LNZzh560+Z/oX/m/Yf/buGUBgYfAgX5jXkG0WyOBn89d9h4/O/zuT//AVURcd5qYvuX/5tIgPtL7t4BgavPN80YgESJneYth//Gdp+/GWXxcDg4vHN8xpiYGDwDWGIhYGBwbkwxMLAwOBcGGJhYGBwLgyxMDAwOBeGWBgYGJwLQywMDAzOhSEWBgYG5+LCiEU5nyFTVF52McgmTyg/xw1mngahKyRSmTOPZZInKM+pmEJXOUmknk/iF5wPWl7+qi49Py8XRiyy8S02j3MvuxgUchlelZCYmpJlYXnrzGNbi3Pkn1swJ51MNo/QSywurDyvTM5AkN7bYD+Vf4F5Pg2C/eV50md2kMqxzKvSeT4CF9burZVz3L0ziSbJ6CYnI0N9bM5NkiiWMFu99Pa0sTA1QUEVYPEwPNDJnetfQ7M4UUpFnE43qqqgYiEavYr1nCHr0icn2GuamLn1dTKqjIzA5q2m73IdE7dvo0pmrM4gHQ12tpN2ui5FyJ7sEs9ZsZcPWY8nMcsgyZZKYB1VoaX7KvUh97nyF0Jn9s57ZBUZUNDNQbRynom7E6jI6LKD4aH+e2eTjG8zu7KDjE6gvp3OpgB3btymrEtUN7XR2lB1nkxZnLpFoqCjS1aGr3aQSKSwa4fcmlxHt9jpams412I8XS0xNzVFQdWweKoZ6Gri9vWvoZqdqKUijnvXRZiJjg6R3l9jefsIoalc7r3K2uwkCUsY/Uof9ZGni4maPdljan4Dk9lEa9cA2b0F9lNFNEWla2AEnznDV9+exutzUS4p9I2MUTxYZXUviSzB5Z5BLKVD5lZ3QVdo6hqi1mdi6u4EJV3C5Q2wMTuJL1mgr7efk805DtMlFE3i6kAXd6cm8aWKXLncwNZegYGeZoSaZmrhiLZ6OxMz65jMVnqHruKxvXq35qtXonOytTRHoKWXtmoPe4t3WYulKSYPCHW/QWvIweHGDFKgldFLYZYnr7OXKHCcVfi2T0dRUzu8PX3Id7w5xtr0DQ7TCvV+67nyLeVzaEIinU7TMfZpwi4zd6+/xVHCRUqx8Oa1KCZJInu0SrFUaV5NVSiWZeR8Cl9DF72NPr7051/ize/6LkzFE+4s71If6jxX/uXjNVLmel4fbiJ/sMTXVxV2V+bwNvRwud5PbHmS1f3E/fNn51cZfuNbsMvw3te+Sr52lN3DNJ/5m9+J+dz7rGjEjjKMXPskLpsZoeXI5wtUX7lEU0ymu63hnOmAbLbROxQFBDe+fh1NNHGSLfMtn3oTLbvP1yZifMebY2zO3uQgkWNjPc7rn3gNrZDgvZlVmptaqA63nVtc30cwPbPE4OufxGmWUbMHzGcsvDE+iF5K87Wbs7w2UINwhBgdHSBzsMbaVgyROOBS9zB1ARcguP61DYZfv4ZFKvPW23egxoGztpPBhkooRi19SMvVIZz5PeYKTl4bGyCzPcViTKGhsYlLV6/iVg/JF0r32zaXL6GVNcrWAN821vOU9XpxXFixyOcVqj1OkCQCAS+7iQIOs5OQzw5A5uiY7WyGwtE6SHY67CZ8Xg8mGXTZjC9Q6WxmswldffoQaTa7E6e9Ei/T7bSimb2MdNdz8/rXcQRqaQ0/cPK9DWkkKwGPDQkJj9+LRQJkEzxFiLb8SRJPpBsJsHlDOEwx8vkygcZKfXx+L9uHBSrhcjR0yYbtXphBh5WyohMKh55CKADJxPj4ELNTtylhZ2ig7fy/fYT0wRaTy7s4bBb2DlMMAl63G5MMQrY8dF2UUpGj3R1u37oFQHVVI5TiHy1joaPoFhynQYxK2Rwunx8JMNncmNQCAomQ34skgWy2ousKg9FRFufmWJ8v093fz9HeLpN3KuWpqmsgm9rGX+t5LLtCMkE8dsCtm0lA0NBq5eDorHKJyj4hkonqsOuj1e0FcWHmLKCy+Yo43QMkEHQTix2i6xrbu4dEwpULdi+wjb+mmkCgiuHhEQYHruBxWE5TkR5K8aOWpJBLc5TMo2sqx+kiLocJm6eK0bExCodblGU7xXwaXdc52tt5YLLxG4uc4a6KkNzdQdd1UvFdijoEQl5i+3F0XWd374BQ+F7nNWE3KyRyJTSlSCKn4LCZnroMQgiEycHgcBQ/GQ6ypdNWkNFUpXL8nGnFtrdo7BlioLcLq3T6K0nirOsim20EImF6+gcZHhqipSGCWZYolTWE0IkfxNHPO2koyThMJY4yRXRdw+r1kz3aR1E18okYOP1ntoqiQUfvID2XQqysxwlXh2nv6WdkeJi25loCQS97ezF0XUdVNUySoKzqOEMRfB4vg0PDDF29SiTgwiQJFFVHMtlQSlk0XScR26Go3avDqx1VxfS93/u9P3n58uWnHdO9cHRNYX11hXgsxl4swaXOLvKHW6xubGMJ1NFWH0ZVFdz+IBYJ7O4AejbGytoGx5kCwVAIXVUJBAIgdDTMBLxuNFXB6vLhsJ5v1y9VKePyh0jGdymXC+xs71LT0k3ArjMzOc3ufpxA7SXqa2ooJXZZ3doFu5eqUAiHTcbm9uGwmCgrCoFgAAmBqksEfI8/nc7CZPchFw5YXtuibPLSUOWjpqGJ3NE2q+tbmHw1tDdUoSkK7kCImrCPlYV5dvYPuNTdj99pRVE1ggH/+RtfKCzNzrCxtQuuEG31VaiqIBiMUEjuEEuWiYQCTwx5+CBur5v1hTmOUgVq6uoIhvyo5cp1kYSOJkyV66IpWF0Bmqq9zM8vsheLY3H5qAr52FxepKxLrK+u09zUeM5tKyXC4QBriwts7+7jCjdS5dKZX1rmKF2mv78biyzQseDzOhG6hpAt5A63WVrdIJkXdHe1U18dZGVhgZ29GLLdTU1tHfnjStsXhZXGGj9L84s4w81UOVUWlleJHR7jC1cTcFtYnFvC7q/DI2VYWt2kKNmJBIL4vU4w2fG47Oe/Li+Q1dXV3DdNWL1nzZ3rb9M9dg3HhRqbfXxQCgn2E9BUF/jwkw2+Yb74xS/GL+ycxcumoaWVM3YkMHhBWBwBmhwvuxTfXBhi8RGpqq172UUwMHihGINoAwODc/HxEAuhkUpn0dUSmVzxzFNy6RTqh9i0y4UchbL6TIqknZalVMg+szTvUS7mPzTNQib9kWzpQgjS6dRztyZn0unzf8l4AWTSKbRzlOesPpLPpFF0QSaderhOQieVPtuOfxH5mIhFiZm5ZXS1SCpTOPOUbCrxoWslSoUM+dKzubFL2QOW1vYp5ippHq7Oc1J+NjdHYn+D3UT2A8/ZWZol+ZEWhwgSiSTPb3O+CovzM5QfyaScS7KxHXvOOZ9NOpk4l43/rD6ytVhp62QigfZgGkJlZm7xnCUQz7SPPA8uzJyFmk8xObuIpqkEGzpoqw+xsTDJfqqISRaUNRu6XiabUzjaPWFhPYbFYkbRTYxEh8imkrjrmpm7+x7pMgjJwWi0j52lafYSBcx2L00hK5rLzdrsBPFcEVkIhMXH6NVudlZmOcyUiW2uUdc7ykB7I/IDn+zyqQOm5lZB6FS39lB9+gWslM9S1q3MT01iPspxpesKVb5HZuaEIL61zOreCRLQ0XsVc+GA+bVddE3lUs8QVS7B3dsTaLKZQipJ/UD9Y22k5E947/YsFquFVPyIwV5IH24zvbSNjE6woYOOpqqHPnEKTWFueoJcWT+1xXeRSaUQao6p5QP6e1oRWo7p+T06m3zcmFzGYpGpauxATu8SyxVBUbDYnCjlMqqq0DUwgt9c4sbtaWSTjNVXzdXuVhKxDebW9rGYZBLp0sOFF4KtlVkmt7KoyNR6BNPz6whdpb6jn7A1x407yzicVlRhwm7SURSFYGMnDV6VG3eWcDjtKBr0Dw3jJM+t21NgMmF2hRju7WBp+japkorDE+FK56WHrl82lSRU38jt6+9QlqygKffba+uMPlLOHXPj9hwWm4XU4QmhPsikklQ3NrO7MsvGYQazDLmShF48ZHZToa+zDrV4wsJGloagYHJ+C7vdSlmVGBrqY+K0j/R19xH22r7RW+aZc2HEwuz0MTQSBV3h3VtTNPt1dtJmro2Po2b2+PLtHYSmkMuX8Ik0llALY931JLZmWdg8wpzNogmN+HGe17/lTWxmGSW9y1bayrXxfiRgf3WWklWjkD4i0nGN9pCN6XffJqUItveTvPbGNTJ+2LaFH+poIJidXqRv/BM4TRpvffVdqgZbACgXCyg2M/X1jUQGh4lYz/6EsrcXo70nSpXPgRCC63fXGfnEG5hFga99fYpyxIK/uZf2Oh/Lt//6jCGzYObuNFei1wjYZN798n8EYHp2heFr34LdBO9+7asU6sI4Le8PKBN7y6juJqLt1axPvcv2cYFsNocQGtnc6Sjt9N+ZeAZnXQdDrWEkSWJhZ5Lw5U/QFpD5s//4Fb7zv/gu9OQu09txTIkNeqJv4LdKzN94i71sExuLm0TfeBObLPjLP/+Th4svSdQ2NZOx6rQ3Rrjx9tsMjF/DblJ566vv4e+tB3c1Y9FObn/1S4R736A5aOWdd25Q21WDZo8wNtZD7nCTmcUNHPk9WgfGqXJZWL75NbYyrRwdxmmNforaM27EXDaLDsSTBT71HW9gpczb707QGlDP6CMq07PTDLz2STxmiXe+VGnrXC6LVs6yEsvzyWvj6IUEf/HOFAiFbP7UyCYUcrkiqkvFHGhkrL+F3aVJ9pOl+30k/IQ+8rK5GGIhBLGtJdb3U5hlnURapZTN4fB6kagIidv2gA1YshAKVAzPHr+H/GoOL4BkYjTay9Tt9xBWHx0BgTtY9ZhvTpLthHw2QMJqNqHoUOU18c57N3FYrPQNPjoy0Dk+iDN39zYAvvBT2lYk6B+OsjA3y0pBp2eg7yFbcbimlnx6l2Cj67ROYTKPFlpAXjPhscqnFvgw9+3e5srJboeNUll/SCwyh0fspFKUE1sILFy2y5z1IiCAUNsAudUFrn99mcbLPSDbCHqtSOh4Qz7MkoRqNqNrZUqqCa+tkk8k6CaWLKBLVqymilszEAw9uT2EznE8xszdSv0D1XUgyQR9lfo7XS4cDhtIErIESDKhQMXU5nC7UYu75FQZn90CkkR1xM3KcQGH04vP9cFrgAI+b2WhHzKSBIVE8ow+IijoZtyn7Vhp6wpqqYjNUdn1XrY58Tof2af2nttVMhEJVOpjMVvI6M9tifAz48LMWWxu79N7dZi+7nbQNWweD/nkMZouKCQPyZYeiHUhFHb3T9CFIL5/hD986lYUArPDz3B0DFsuTtEbIrm/g6LpaJrGg/Zv6ZHuoeoyrW3tdFxuxSQ98lSXZMKRIM2dfYyMDHOl69JjAmSWoaRoCF3l4OjkoWNCgIaJ7v4hei4FWd04IFQdoaN3gJHhYTpaG/B4nRwfJRBC5zi+//C7caXAeKyCo2wRXVM5OIgDJuwmhVS+jKaWSOZKp3bv9/FVVxMMRBgeHmHoaj8+l+20Sha0ch5NF2SO42SLZTRNo761m+hQN6vLq6etJN0vgPRAYYIuif1kAV1T2Y6nqQ67MFMiV1LR1BJHR48vlJAkCVVVEciEIiFau/sZGRmm+3LTB3dUobG7f4iuC04OD7F7/YTcJvYTWXRdY30vRV31vZv2Q57aj1jPnaEwyf0d1If6iITbqnOcK1fa+vD9B5XZ5qCUT6HqOqVsklQuj2R2oBQz6LpOYn+X0hOs//f7yCs08fsgF8PuLYHHbmZ+YZFUXqOmpppwVQ0OkWVheY102UxDVQif14UqzJj1IulshoP9PYomH92tdajlMm6/h4WJu2zt7mPyVdPa1IRLzrGwtMphMk844MXicGOVdFz+EBYZ1HIJu9PK7s4BilIilTxideuQxrqaB979JcKRIKsLc+zs7VOWbATcdjQseBwWzE431SEPizNzCF1hbS9JU93DS8N31hZYWt0gkdPo7GynvsrH4vwCu/sxsLmpr6vleHeVje19bO4QkUgYp83yUCOFq8Kszc+yGzskGKomEKmiLuJlaX6O3b04TZ39BNy2h7qozR1Ay8RYXtvkKJklGA6jKWWCoSqsWobFlXUyikQ4GMaiZZmeWyR+mKC1oxO7CZz+IFYJiqUy4VAQhIYqzLS3t7CxMMPW7j7+hss0hDwEfE4W5hc5ODqhtq6JYDCA6YHXOZPZxvHuGqmSRNflZpYX5tjd20c1O/A5bQjJhtftQCmXcPqC2EwSpVIJt9PM4eEJJ0dx0qqV3q5Wqqqr2V2dZ3N7F3dtK80RH0q5hC8QwnSGXpTLJXyBIGq5TDAYRAKKZYVITQNO6fE+0tJYw9LsDPvxQ0LhWgKRCChlApEa/FaNucUVkjmVuupqQuFqtGyclY0dinLF3u1125CtDtwOG5qqINtc1Ea8LM7MYXb58TjOtwr6RfGxtXvvr85SdDdwqdr3TNIrJ9a4vqzyRvQypewJN6fWufb6COcMgfEQmZM4BclNVeDVXmF4kcgeb7J2bKK/4/xL5Q2ejo+t3dsTqsZpeXYLciz+Fi5XrzFx9y5Wh4do9OpHEgoAT7Ca8y0ZMzgvVqefWunCvFFfWD6WYuH2hz/8pKdAkmTqmtupa36myRo8I6wOHxFjnchzx5BjAwODc/GxFQshdDKZs12OuUzm8a8JLxuhkcmcHZC4mM9S1p63p/LFU7kOgkwm83y+AAid9AN9QOgqmeyzCfYrdIVM7my38EdPVJDNZF4pG/yDXGCxEMRXF58cLVkoTM3MnXloeXaSwgu494QQbC0vUjqHMglRZGp2+cxj+2uLHOfKz7p4LxUhBEuzk5R0wfHx8UeOWfbBmZSYmJp//3/LKabmVxF6mZWl1W8saa3I8YdY7j9CqszNzrx6D7JTLsycxd7GEo5ICwGXlZ3leexVddyeuIPnOEtv7wAB55OqIliZnSCRV8HqZri/C6EpzNy9CaqK3VvNQPclTvbWWdiKg67T0tVPnV/i9s05VKHTdLkbr5xnZmkToam09Y0Q8dof+2IvhGB1boLjnAJmFwOd9dy4fZuGTIm+K1dwPeJxEEKwtTjFXrKAySyh6laErjI3eYdsWUeTbAwPD94/v5w74fbEPJIMvppWulqqWZy+SypfxlfVSEdjgNu3p9CBQG0rl5urHy+jXubOjZuosgVF0fB7HJXgsTYPwwPd7K/Os5/IoWFhaGiA0skuc5txSskDFHsVb4x1cOOdu5gdNpRiiZ6R1/FbFGamZyirKq5IM92tdWe4GXSWpu6SKmlg8zHS13H/+uRzlRHV1tIUO8d5zBYzZpuHKy1eNo8tdLSEKaTj7KdkmkLWU9u/Rqixg9b60FMHozvcXuLG3WXKspXu9sbH20grMXV3kpKu4/DX0ttew813b6LLFnS1TFPXIHU+jXy+ROpwm5mlbcxmGdlsR9ZLlMtl6i4P0FTlPaP9NeYn75BTdCyeKga6WkjFt5hd3cVslkm+wg+FCzOyKObeH4oXMmk0i5OGhib6rw59gFAASLT1DDIyMoK1lCSn6JSVEvXt/YyPv4Ylt8t+Isf0yj7j4+O8NjbM0vQUCJXtwyzR8THqwl6mZ5cZio4xPh5lfmLizPCd5cQ6xyLMaDRKgzPHRspCU3MTAwN9jwkFgJaNs5U2Mz4+zmBHPTlFI7W3RMnVxOjYOFcaPcwsbd8/f+L2JL3R1xgff53i3iInRY3N7T2uDI3Sdamemdt3aR2IMjo2Smx9kbMXnersJYpEo6P0tgQ5LDkZHRvDpaXJFDUa2nuIRqPUeQUHyQJzi+sMDQ8zPjqM2+XGgspxQWJsdIxr4z3Mzy5jsjroHxohOjZOJrbxhHxlLvcNMTISxZQ/pvzAbZROpVFzR2ycSLz22jhXO+uIHZ2gq0UyuYpNWlNK5Aql+7b/aHSIg+3VpwyjWsmzqqGRxqY2es4QCoCtpVl8Td1Eo2OUjrZIF8rEEiVGx8Z4bXyQ9eUV0BXSmTxKMYPsq2dsbJzS8T4NXVcZf22c3ZWzF5BJsomeq1FGoqMoiT0UYGZhnej4a4xGh9GL6aep0AvlwowsHuT84WFBLaa4dXcOk9nC7nac5n6B1ebC566YXnxeB9l0BovNhSxJSGYbFnR0oCoSxiRJCKFytLd3334dqKo+M69s/ID9mM6tQgyhC5qqJT7o0pcyWZz+SqBYi8uP23pELpHBX9eOBDi9Acq7cbAD6JR0K27rqcXY6ySTVfAFgthPbceJkxMK03eRJbC6fE9spaDfiyyByWTBH3AAArPZhFYqcGd6Bk2ykDzcpyNwmfbmCH/91XcIeey0tHUBZcJBP5IEwmwDvUz6cJuZlV2sFjPx4ww68Kg0qvkENybmsVqtbG0f0DX6QOkkKGezOH2+B+z7j67fqFz1w+1lVvYSmCXBSbp06qd8EtLDbVwG8ZkAABklSURBVCDE4397DEHq6IiTE4XDTRnV5MJikggF/ZXP5bIF6cE1uZKJoM8JQuDyebBbzSCJJ+ZSSh9wa3oFm83KTuyEPqEhJCsWkwTCRCAQ/MDSvUwujFhYzSZyxRK628JhLIa3k0q0ZE0gzDwxaGtibwtH7WX6Gv1kDyqrHsrFHMeJPJ6QnaOTPHVX/MS3VikrGrKWoyybkXk/TUkyEawK09k3iMdmQtPFmcFpPTU1BDJFhoY7QWhIsoltIdB1gZAfL6PN6yG3FUfX6ygmj8iVVbxVIRb292gJNpE4iuP0+aFUAGQ8No3jbImgw8RBMk9Hh5WK0VgCSRAK+vC199AQcKJpGuYn3kVnH8inDilaQ7zW38bU9SQCEMUSde3dNAds2Gx2EOXHrPBb6+u09r1G2FrmYP+tM9M+2l7D29JLT7Wd5P7+w2UQYPV4yK/voOuNFFNHpIslZLONcjGDEDqJ+B6K3Mja5i590TewqCn+01sTgE6hqGC32x6vlWTFquZI5sv4HGYOYzFcXj8SMrp2aquWHq2NRCASwuxoorspjKZpmKQyHxSNWEL6wOMPsr+2TKRzmDa/xNFeDDAhU6KoaFgpc3xy8qFpvCwuht0bcHk9rM/PsrsfR7Z5qK2vw+8yMT+7iMMbxmV/RPeEoFAs09DUxM7yPPsHR7gDEaqqI5iQyZ7E2NrawV19iaYaPwGniem5Rfbjx3Re6cdlkykUdcIhHyARDriZm51jbz+GbnHidz/+YV+2+yC3z/LaFvGjE/zhapxymcWVLXzBCDbLw89b2erCVDphcXWTZFGiPhKgur6JwvEWK+tbZBQrfd2taOUiNo+fhtowi9PT7OztEW7qpDbgolAoEgxVVsGGq6tYn59mezdGqqhTFTojgrfQKRQr1mxdLaPKNgJuB+ViAV+klvzBJlt7cWyeEKGgj8PDONlkksTJEXNLG7S0NFAsCcIhHxI6+YJGc0MVi3NzHJ1kCdfUEAkHHzOtOTweNhdmiB2c4AlEqKqpQink8YXCKMUi4ZoGrEqKhZUNErkiQjfR1tpO9nCD9e09CsJKJBymNuhkbmGZRKZIVXUNIZ+VuzMr1Nc+Pj+DJFEV9jI/PcPu/j4FnFzpuoRJtpA73iaWKlEVDj52n3sDYQ43l9jY3uU4WyIS8lMqKoRDARCCfLFMKOilWJbwu61IZgcep41iIY83EMYiQ6FQJBQOPlYml9fN6sw0B8dJ/OFqItURgi4Lc3NLHBwliFTVEY4EH1nV/PL52Nq9DZ4NejnHW1+/y7VPfgLUAu+8c5PXv+XN5x+oWM/zzo1FPjF+9TlnZHBePrZ2b4Nng2Rx0tfVxNTEHWSzjZ6rwy8morlkobHeeH69ahhiYfBEJEkiVNNEqKbpBWdsoamx9sXmafChXJhPpwYGBi+Xj4VYlIt5yurjkYaEEOSy2RcSTCSfy54rOvSzpJDLfmjE8hfNi2qHp6m70BWyT4j6/g3lLyCfzT7BV/Lx42MhFtnkEZknROU+iMd4EQHLjuOxx6JVP28SBzGKzyVPQSFxwP5x6il/JlianaL4Aho8cRCjpMPe2vIDGws/VJj7x4RWIHaYfKb5r89MkNUEC9MTD0S++nhzYeYsDrZX2YgdITQdu8tDOZ9D0VTaeq4ilRVkIVifn+IoV0RXNSyeKq72tFIulUAvc+fWbVTJTFkVBD02svkSZleQwSvtD32mUgopVndTdLU3oRXTLG0nqfUKFjbiCF3QPTBE8XCDzfgxkgDN5GJsuLeSjwQH2ytsxhKoGgyMjJCPb7CyE0dCYLW70UoFFFWhuWuQuuDZAXCEEKzM3OYop2G2WnB7QlS5BWVrmNqQm6PddXRPNcppniszdzjKKQjJzshIP5ZHvluuzU1ylC8hVA2rt4bB7orFeG59D3RBc1cftR6Z23em0CUJT7AOJT7PdsFGX18/paNNUvkyrkAtHrmAt74Vn93C9tIc/rYe5HSMybk1TGYT6XSBy2fVSS1w984kigB/dTONPsFmUqpY1mdnae2+QmJnhY1YEh0zg0MDxNeXSOZzCNlF35UOVucmSeZVXMEaXFoJpZDm3Zs3qU3k6bvSw87CBJlyxUZ9pSlw/1hvZyPlkoLQysxMTpBXdCSrl6GBbnaX5zjI5tFVDckeIDrQ+djnzkR8k6I5RG3Izcn+JmX7vRAI984UxDaW2T5MowmZweGrJHdW2To4Rtd0HC4PpXwOVdNov3KViFti8u4kJQ3C9a1U2cvMLG+B0Klr66Wp2vdK7qd+YUYWxcwxllAro2Oj7K2t0zU4QnSgm421TYq5DEVFJ30cI3Spj9GxcaTUHhkVUskEQmjsHBcYjkbprndxUHIRHR1Fyh1WQuA/gNnm4uRgD13Awe4mFoedmeU9RqJRhq60MDu7SCF9iDl4iejoGCEpw1FRI5Oq7BkRqW9lZGSE7kYnq9sJitkTZF8jo6NjnOxscunKINGrvWyurDzRSagkN4mVA4yPjdJVa2f7KEspn6FwOnoq5bMUyxrZVAJVaOwcpLk6PMLYSN+ZRqzkUYyq1n5Gx8YRyR2yisbkwibR0THGR6+yND1J9iSO4qwmOjpGd3sjdU0tXO7qpbkmyObWFm29V+lubySXTqGcPslzqRSqEMxMLzAwOs7o6AiUzvKsCpamJqnrusroaJSDzWVs/hq0ow0W5qdR7CFM5QTLsSKjo1GuNDiZXY2Rim9hr+lksK+LTGyZvLWmcry9kVwygeTw0djUzMBgPy6bmY7+YUaio5QTewin//1jFo1kKsf+2hxy4BKjo2M0uMos756QPdnD3dDD6OgYjvwBqTP2WikXsu+3/RM2oqpuamdkZJjWKjObe2kK6UMsoVbGxqLsra3TOxRlpO8yGxvbrExPEmjuYXR0lNb6MJMzSwxGxxgfG2VrfuJ++75qXJiRBZKFSMCJhIQvHMRulpExg3j/ZjeZnYR8diRJwmYxoTzwMhkK+DBJEhazDX/IhySB2WxCf+SFU5JNtIYsbBznOT7I0NPfyMz1Xe7evgUI/P5aKJWoDrmRJAm71ULp/spXwdzkTXKqiXLmAFdDGCQLYb8LCQlP0I/DakEWysOW4UfIHR7hq+1GkiQcgWqcj2y88/AcjImr/R1M3b6ByRlioPfyY1Zrs9VF0GtDkirRystqGZPFhdkkI5ns2CSBPdJEY26Z965fp6algwfHPF5/ELfdcoZLVgA6ZWHBaZGRgFA48niFBJwcHXOiTLEtg2xzI5BpbWvkC3/5Hj/w/f0UD9c5jO9x61YJhEawNkwh6aImXGnnzHGSQGPrE526av6EmxOLWG1WdvaP6T/jfsumCwQu+5EkiWAoyM5+DrfsoDroPL2WJsqa4AO/D58xHyM0lZmp2xR1M7lknEh7PVbJetpfZXzhSrxQzBaEppEuKHR6XZW6CBVdsmE3y0hIuG1mFFXHanp8LdHL5sKMLCpDvscv4mNBrp/ofDvvwE6iuq2L/el3EK4aHDY7vlCY/qtDjIyM0NVWf/+8x8qi5YlnTERHhmiq8t2f+LpnKH7UWFzKpckWlUeTwRUOko7FKxO0xzHyOljMZoqlEkLonBw8PA/j8lczMjqGJbPHYeHxCQOJh9tFki2gVSaF1XKeEjIyEnUtnYyNjbC1PI9AQtV0hBCn5a783maWyJcUhK5xdBAHZKySQr6soesqx8ePR+1GgkDQR317DyMjI4xHBzAJlYWlLT59bYDJ2VVsXi++QIih4RGGR0a5VB96qM08QR9H+5U20fV7QltZg6Hpgv2VBYKdwwxd7b8fov/esXv4Am6OD48RQnB4eIQ3UDEuP7nPVDCbLQ+0/f4DbV9JWykkSShORkaGqA95HngMnJ2u12niIFGJ4aELGYtUrrSfqpApqVjMr+ZteWHs3uVSHqvLh9NqJpfLEQqHkdEpFDU8LgtWlw9JLeEJRrDIUMzncAVCaMU8gVCIYqFMOBxEU0qoJgcBt41iPo8nEMRieuTiSBZSB3GaOjtx2W0VK/jsIvuxGLLDi03Wsbn9OK1mysU8Fk8QqVzAG6lFTeywvh0Du4eAN4DTKjA5PLjtFvL5HIFQGJOkky8oJPdX0d3VeB2Wh7I3OfyUTzZY3dwlWVAwS1YuX77E7uo823sxypKNmtpaZLWMy+9l9s4ttnf3UWwBLjdWP2YVLuZyeEIRLBIU8jk8oSqq3CamZxfY2z+gvacfUznJnYlp9mMxwvWt1FeH2FheoIwNu1kiGI4gS+D1eViemWYvFkdYXNQ1NlLttzMzM0c8fog/VEO4KoL5oXkTiWAkwtrcJDt7+5zkFFzkEZ46murrKCb2cYQb8ZvyzCyuEovFsfvDSGoJdzCCVQa7O0gmtsra5jbpIngcZtzBCC6pxMLSJrXNLWwvzHBwlMATCFNdU4WdyjGP34+uyzS3tnCys8za5g4Fk4ee1gbKhTyu0zxKhRx2fxj7I+G/7Q7Xw21fU4NJU3AHI2iFHMHqegqHm2zuxJAdPkL+IDaTdtpHTORyecKRMJLQKZR02jva2FqaZWtnl7Jkp60hxPTMHLt7e6cR2B8Pf/CyMezeL5m15RWa2toeubEeRi0luDm9x2sjV15gyQwMHsawe79kWi+3f+g5sslOXc2zDUBsYPBRMMTiFUc2O2huMEJXG7x8Xs2ZFAMDg1eOCyMW5VIB5YwI10JXyZ/uUH1eNLVMofT4V4gnIYQgn889FnVZ18rki994zEShq+QLJdRykdIZ3/DPLpNOLv9sIlVfFITQyOWfrW3b4PxcGLGIrS0STz/eUYSSYGJm/anSKueTHD5FZGZJkojv7T4WdVktZogffXDMxPzRPvHkB+elFo+Ymtsknz7hJHPO8PJCZXcv/uHnfZzQskxMnx0B/VVECI2Ntafrm68yF27OopA8YGZ5E03VabvST8gGifg2N26kUVVB79AwHovG9MQkBVVgcQUYuHKZnZVFkvkcuuSirdGPrmmc7K2ztBUHJC73DBDyVrY83Fqa4zCXRyurmFxhhnrb0VQVoSvMTEyQUwQ2d4iuZv/pztoVtOIhqzHoaIlQyh2zc6iQWLtNXHjp7xugsaqy92o+EWd2ZQtN1WnvHcB36r/RdQ1dEmilDLduTyGZraCoXI6Oc7g2z6XOHiwSLC/Mc+lyW6VMWo4b700hmWRUVadrcJig696muoKd1Xn2jrMIk4Phq90szC7QeeUK+YMNklKI5mpv5UytxMzkNAVVwxtupPNSLVvLsxymi2BxMtjXff+rjdAV5qenyJY0/FVNNAbNTM0tI4Qg0tRBa52fmbt3KGoSiqoT9LlIZ3OY7D4Ge9uZm3jCsb5OUvvrLG4dghC09QxQ5bOzNjfBQaaM2SoDdoRWZu40/3u/e7Bsi7PTpAsqnnA9rdVOJqYXEAJCDe20NwSZnbhNXgFdValu6aI5bOPO3Wk0wBdporM5zOzUFHlFwxOqp6u1ntjGAuvxNFarBbPNQ1+b/+FrfaTSXOVkZn4RRVEJN3YQMqf5+o1bJAoqAz2VZQWl1CFTSxvoShHFHubaUPfzvmWeGRdmZHEPuzfM8PAIw33NrK7tAFDExshIlOG+S0xNzbO9NIOj5jKjo6MERZL1gyzJ+Cb26g4G+zoRSp50rsjG5jatPYOMjkYJeN4PEJs53sVZ20V0dAxzeo+UIkgmTijl0xwVTERHR+nrakVXC6TS778KCLVI8nT0oylFUpkCdU0tdPT03RcKAIcvUqnDlQZW13bv/72cz5Irlpi9c5eWvhGiI8OUU/uUdEEqkbhvHkwlTtCFzkkiBUJh97jIUHSUsZEepu5M3D9PzcTYSMiMRKO0+UrMbueoC9qZml1kdv2IuvD7u65uLc3hru8gGo2S3Fshr+g0tHUzPDyMW2RJPBCifn91DjnQTDQapb2piqmJaXquRhkbG+NodYZcWWNz/4Srw8P0XgqzeaQSjY7iUBOc5MpPPHacyjC1Emd0dJTo0BVmJ6dQ0rvs5lyMjo7SVesmrQhi6/Po3kZGR0epsRVY2j6+X7b4xgKKs45oNEpnSy3TdyfpHIwyNjZKYmOWdElnY/eQ3sFhRkcH2VlfIXe0h+KqJTo6RkdLDburczhq2olGo2Ria6TSJyztFRgfHaWvvZad2MHj1zqdx2R30Tc4xEh0hNjGEu5wDY1Nl7h65fJ974vNFyE6MoLXbqHt0sXaD/OCjSwEu2vz7J7kkbUcOVFx+VVFwsiyhNXpA2WNdEanrtmLJElUVwWZSeSwm9+3Dt+jd2CA+fkp1jQzvQP9uG2V5pBkBzVh16kF2FyxAANWV5CuxiTvXb9OsK6FxjNCXD5Y1jMd/kKwszrHXqKArGXJUQ08vKAso8j0uKxIskQkUv3Iz8VjjuNIOIRZlhBWLxaRvx9dO3d0wOFhgtu3MqArRJohUNXMnZu/T+3w38J833wkSBwckE4oHG1JaCYHqAUmJ2fQMHOwH8PX0nc/v1QqR7jbf9qWOmXdittmRgICHju5gkog4Mcsy5gtNkIRU8VqbjGjqfoTj5VzeWwuHyZZApsbi14md3yCt6YFWZJwhmpwrW+TSeUJXQ4iSRLhSIjd3QwQBgTpRJbQ5S4kSUJCp6Ba8NnNSAhCXgfpnEIwGMRmkZGxIEkCd80larOLvHf9XepbO0nGDzk5LHGyI6PIDrR8Dqc/UOljbj9ex6ObbleudSK+xdJGHLNJ5jhTfOL1T+yvUnDU0OV3fkD/efW4YCMLlcXtBKPREa5cboZT2+/RcQIhBEoxA2YXXo+dRKoSx+LwKInf73zM8gxgcXjpH4rS1xZkbnHroWOPWrMrf5Sobmxj/LVxkluL5B5xVstmG6pSqNi0Tw4oV4JHo+nigfUcKku7SUajI/S0NSLE45O2DpNGplyJPn1yclhJG3G61kUjcXL80PmHxwl0IRBqljLO+xfVGQjiD1QxMjLCyOhrNFd7OdpZJdJ1jcTGHGX1Xt4SnoCPhrYuRkZGeH18BCW5j/A1MjIyTJXX/lDHd7tsnCTSp3WSsZlU8oqOEDrJbBGnw/yEdST3mvHsYyabnXL+1Aat5FFkC06/l+xxxaJdSh2R18Djc5I8SSKEIHGSwOW9Z0CWcHvsnBxVjglkHGb1tC0hkS7gcd1b4/JAGSQTzZd7GB8bZm1xDlfAR/2lzvtt4fO5KWQq9VXzaTKF4pnXemV1k+6rIwxd7cOkKYBUuS7i/euva0Xm1g7p7Wg6b0DwV4YLM7Kwuz3IFhsd9T7efe8GTtepWUm2Uh90cPvWLRRNMHB1GLdZZeruBDe2BGZngMFqD9vJwP3Kmq1OPE4zq3MTHKZLCCHoGhi+n5fbH7i/etPlC2CVJXz+AGo+we2JOUwWM7ZwEx6bHZ/nfcWQbGF8rHHjxk0kE0QiTiIRP+t359igk0v1YZDMtNd4ePe9G7hcDuqrwsgmG36fC6tDxyVbaRse5OadG5gsFvJqxQre3trE5I13MZlkfDXNyJJMwF+Zb3BIRW7dvIWqqAyOjNzvhBZ/A23Bad597wYmWaajr494WtB75RLFiJmNvSM6m6oAaO0ZZOLuXW5smrC6A/S216Nv3uVmcg+zrwan5f3nSkNHH9MTd7mxC/7qJvoHrzBx812QIHypF7fVRMBfGXaZrHZ8bg2QcHp82CzmJx6zO1z0tUW4/u57IARXBgaw+hxU797lxs0jLDYHHfV+appqOZma4EZ8DdnuYbDvfdNabdsVTiYnuHFjDW+4gf6r/dy59R7IEGzuwWeT8Z/u1QISAb+f7Mk+UwsbmEwStc1tXGoIVuq3I2Nx+envvkxreJ/3btzEbJFw2GxnXutguJGZ2zew2Rw0tl5CkqzUeiRuTswzNNCNWYL4xhJ5DSbv3MYTrqXrUsMzuT9eBIbd+xVn+fZ1PFfGqLGfPQgUapLrt3d4faz3BZfsmxS9yDs35vjE+NDLLskLxbB7XwAC1bXYnrxbEEg26moNO/gLQzJRV1v1skvxUjDE4hUn3NDygcclk4OWJsMO/sKQLFxqvjivDs+SCzbBaWBg8LIwxMLAwOBcGGJhYGBwLgyxMDAwOBeGWBgYGJwLQywMDAzOhSEWBgYG58IQCwMDg3NhiIWBgcG5MMTCwMDgXBhiYWBgcC4MsTAwMDgXhlgYGBicC0MsDAwMzoUhFgYGBufCEAsDA4NzYYiFgYHBuTDEwsDA4FwYYmFgYHAuDLEwMDA4F4ZYGBgYnAtDLAwMDM6FIRYGBgbnwhALAwODc2GIhYGBwbkwxMLAwOBcGGJhYGBwLgyxMDAwOBeGWBgYGJwLQywMDAzOhSEWBgYG58IQCwMDg3NhiIWBgcG5MMTCwMDgXBhiYWBgcC4MsTAwMDgXhlgYGBicC0MsDAwMzoUhFgYGBufCEAsDA4NzYYiFgYHBuTDEwsDA4FwYYmFgYHAuDLEwMDA4F4ZYGBgYnAtDLAwMDM7F/99OHdsgEAMBEPS9qMA5nSICCrTkHtCHdglHAwSX/QczFWy0ZgGUmAVQYhZAiVkAJWYBlJgFUGIWQIlZACVHay2vjgBuL4+995npF8B/mdnWWudjzvmKiE/v/RkRcXUYcB+ZmXvv7xjj/QO2+QQ+H0iWvgAAAABJRU5ErkJggg=="},{"background-color":"#383E41", "background-pattern":"" , "items": [], "preview": "iVBORw0KGgoAAAANSUhEUgAAAQsAAACWCAYAAADJ2q17AAAABmJLR0QA/wD/AP+gvaeTAAAAsklEQVR4nO3BMQEAAADCoPVPbQwfoAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA+BtyfAABMgdIAQAAAABJRU5ErkJggg=="}]}